library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.ReSamplerTypes.all;

package inputs_test is

-- Declare constants

  constant inputs :inputarray := 
  (
("00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010000", "00000111", "11111101", "11110100", "11101011", "11100011", "11011011", "11010101", "11001111", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11010000", "11010101", "11011100", "11100100", "11101100", "11110101", "11111110", "00001000", "00010001", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110110", "00110011", "00101101", "00100111", "00100000", "00011000", "00001111", "00000110", "11111101", "11110011", "11101011", "11100010", "11011011", "11010100", "11001111", "11001011", "11001000", "11000110", "11000111", "11001000", "11001100", "11010000", "11010110", "11011101", "11100100", "11101101", "11110110", "11111111", "00001000", "00010001", "00011010", "00100010", "00101001", "00101111", "00110100", "00110111", "00111001", "00111010", "00111001", "00110110", "00110010", "00101101", "00100111", "00011111", "00010111", "00001110", "00000101", "11111100", "11110011", "11101010", "11100010", "11011010", "11010100", "11001110", "11001010", "11001000", "11000110", "11000111", "11001001", "11001100", "11010001", "11010110", "11011101", "11100101", "11101110", "11110111", "00000000", "00001001", "00010010", "00011011", "00100011", "00101010", "00101111", "00110100", "00110111", "00111001", "00111010", "00111000", "00110110", "00110010", "00101100", "00100110", "00011110", "00010110", "00001101", "00000100", "11111011", "11110010", "11101001", "11100001", "11011001", "11010011", "11001110", "11001010", "11000111", "11000110", "11000111", "11001001", "11001100", "11010001", "11010111", "11011110", "11100110", "11101111", "11111000", "00000001", "00001010", "00010011", "00011100", "00100011", "00101010", "00110000", "00110100", "00111000", "00111001", "00111010", "00111000", "00110101", "00110001", "00101100", "00100101", "00011110", "00010101", "00001101", "00000011", "11111010", "11110001", "11101000", "11100000", "11011001", "11010011", "11001101", "11001010", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11101111", "11111000", "00000010", "00001011", "00010100", "00011100", "00100100", "00101011", "00110000", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110001", "00101011", "00100101", "00011101", "00010101", "00001100", "00000011", "11111001", "11110000", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11110000", "11111001", "00000011", "00001100", "00010101", "00011101", "00100101", "00101011", "00110001", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110000", "00101011", "00100100", "00011100", "00010100", "00001011", "00000010", "11111000", "11101111", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001010", "11001101", "11010011", "11011001", "11100000", "11101000", "11110001", "11111010", "00000011", "00001101", "00010101", "00011110", "00100101", "00101100", "00110001", "00110101", "00111000", "00111010", "00111001", "00111000", "00110100", "00110000", "00101010", "00100011", "00011100", "00010011", "00001010", "00000001", "11111000", "11101111", "11100110", "11011110", "11010111", "11010001", "11001100", "11001001", "11000111", "11000110", "11000111", "11001010", "11001110", "11010011", "11011001", "11100001", "11101001", "11110010", "11111011", "00000100", "00001101", "00010110", "00011110", "00100110", "00101100", "00110010", "00110110", "00111000", "00111010", "00111001", "00110111", "00110100", "00101111", "00101010", "00100011", "00011011", "00010010", "00001001", "00000000", "11110111", "11101110", "11100101", "11011101", "11010110", "11010001", "11001100", "11001001", "11000111", "11000110", "11001000", "11001010", "11001110", "11010100", "11011010", "11100010", "11101010", "11110011", "11111100", "00000101", "00001110", "00010111", "00011111", "00100111", "00101101", "00110010", "00110110", "00111001", "00111010", "00111001", "00110111", "00110100", "00101111", "00101001", "00100010", "00011010", "00010001", "00001000", "11111111", "11110110", "11101101", "11100100", "11011101", "11010110", "11010000", "11001100", "11001000", "11000111", "11000110", "11001000", "11001011", "11001111", "11010100", "11011011", "11100010", "11101011", "11110011", "11111101", "00000110", "00001111", "00011000", "00100000", "00100111", "00101101", "00110011", "00110110", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010001", "00001000", "11111110", "11110101", "11101100", "11100100", "11011100", "11010101", "11010000", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11001111", "11010101", "11011011", "11100011", "11101011", "11110100", "11111101", "00000111", "00010000", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010000", "00000111", "11111101", "11110100", "11101011", "11100011", "11011011", "11010101", "11001111", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11010000", "11010101", "11011100", "11100100", "11101100", "11110101", "11111110", "00001000", "00010001", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110110", "00110011", "00101101", "00100111", "00100000", "00011000", "00001111", "00000110", "11111101", "11110011", "11101011", "11100010", "11011011", "11010100", "11001111", "11001011", "11001000", "11000110", "11000111", "11001000", "11001100", "11010000", "11010110", "11011101", "11100100", "11101101", "11110110", "11111111", "00001000", "00010001", "00011010", "00100010", "00101001", "00101111", "00110100", "00110111", "00111001", "00111010", "00111001", "00110110", "00110010", "00101101", "00100111", "00011111", "00010111", "00001110", "00000101", "11111100", "11110011", "11101010", "11100010", "11011010", "11010100", "11001110", "11001010", "11001000", "11000110", "11000111", "11001001", "11001100", "11010001", "11010110", "11011101", "11100101", "11101110", "11110111", "00000000", "00001001", "00010010", "00011011", "00100011", "00101010", "00101111", "00110100", "00110111", "00111001", "00111010", "00111000", "00110110", "00110010", "00101100", "00100110", "00011110", "00010110", "00001101", "00000100", "11111011", "11110010", "11101001", "11100001", "11011001", "11010011", "11001110", "11001010", "11000111", "11000110", "11000111", "11001001", "11001100", "11010001", "11010111", "11011110", "11100110", "11101111", "11111000", "00000001", "00001010", "00010011", "00011100", "00100011", "00101010", "00110000", "00110100", "00111000", "00111001", "00111010", "00111000", "00110101", "00110001", "00101100", "00100101", "00011110", "00010101", "00001101", "00000011", "11111010", "11110001", "11101000", "11100000", "11011001", "11010011", "11001101", "11001010", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11101111", "11111000", "00000010", "00001011", "00010100", "00011100", "00100100", "00101011", "00110000", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110001", "00101011", "00100101", "00011101", "00010101", "00001100", "00000011", "11111001", "11110000", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11110000", "11111001", "00000011", "00001100", "00010101", "00011101", "00100101", "00101011", "00110001", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110000", "00101011", "00100100", "00011100", "00010100", "00001011", "00000010", "11111000", "11101111", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001010", "11001101", "11010011", "11011001", "11100000", "11101000", "11110001", "11111010", "00000011", "00001101", "00010101", "00011110", "00100101", "00101100", "00110001", "00110101", "00111000", "00111010", "00111001", "00111000", "00110100", "00110000", "00101010", "00100011", "00011100", "00010011", "00001010", "00000001", "11111000", "11101111", "11100110", "11011110", "11010111", "11010001", "11001100", "11001001", "11000111", "11000110", "11000111", "11001010", "11001110", "11010011", "11011001", "11100001", "11101001", "11110010", "11111011", "00000100", "00001101", "00010110", "00011110", "00100110", "00101100", "00110010", "00110110", "00111000", "00111010", "00111001", "00110111", "00110100", "00101111", "00101010", "00100011", "00011011", "00010010", "00001001", "00000000", "11110111", "11101110", "11100101", "11011101", "11010110", "11010001", "11001100", "11001001", "11000111", "11000110", "11001000", "11001010", "11001110", "11010100", "11011010", "11100010", "11101010", "11110011", "11111100", "00000101", "00001110", "00010111", "00011111", "00100111", "00101101", "00110010", "00110110", "00111001", "00111010", "00111001", "00110111", "00110100", "00101111", "00101001", "00100010", "00011010", "00010001", "00001000", "11111111", "11110110", "11101101", "11100100", "11011101", "11010110", "11010000", "11001100", "11001000", "11000111", "11000110", "11001000", "11001011", "11001111", "11010100", "11011011", "11100010", "11101011", "11110011", "11111101", "00000110", "00001111", "00011000", "00100000", "00100111", "00101101", "00110011", "00110110", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010001", "00001000", "11111110", "11110101", "11101100", "11100100", "11011100", "11010101", "11010000", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11001111", "11010101", "11011011", "11100011", "11101011", "11110100", "11111101", "00000111", "00010000", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010000", "00000111", "11111101", "11110100", "11101011", "11100011", "11011011", "11010101", "11001111", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11010000", "11010101", "11011100", "11100100", "11101100", "11110101", "11111110", "00001000", "00010001", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110110", "00110011", "00101101", "00100111", "00100000", "00011000", "00001111", "00000110", "11111101", "11110011", "11101011", "11100010", "11011011", "11010100", "11001111", "11001011", "11001000", "11000110", "11000111", "11001000", "11001100", "11010000", "11010110", "11011101", "11100100", "11101101", "11110110", "11111111", "00001000", "00010001", "00011010", "00100010", "00101001", "00101111", "00110100", "00110111", "00111001", "00111010", "00111001", "00110110", "00110010", "00101101", "00100111", "00011111", "00010111", "00001110", "00000101", "11111100", "11110011", "11101010", "11100010", "11011010", "11010100", "11001110", "11001010", "11001000", "11000110", "11000111", "11001001", "11001100", "11010001", "11010110", "11011101", "11100101", "11101110", "11110111", "00000000", "00001001", "00010010", "00011011", "00100011", "00101010", "00101111", "00110100", "00110111", "00111001", "00111010", "00111000", "00110110", "00110010", "00101100", "00100110", "00011110", "00010110", "00001101", "00000100", "11111011", "11110010", "11101001", "11100001", "11011001", "11010011", "11001110", "11001010", "11000111", "11000110", "11000111", "11001001", "11001100", "11010001", "11010111", "11011110", "11100110", "11101111", "11111000", "00000001", "00001010", "00010011", "00011100", "00100011", "00101010", "00110000", "00110100", "00111000", "00111001", "00111010", "00111000", "00110101", "00110001", "00101100", "00100101", "00011110", "00010101", "00001101", "00000011", "11111010", "11110001", "11101000", "11100000", "11011001", "11010011", "11001101", "11001010", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11101111", "11111000", "00000010", "00001011", "00010100", "00011100", "00100100", "00101011", "00110000", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110001", "00101011", "00100101", "00011101", "00010101", "00001100", "00000011", "11111001", "11110000", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11110000", "11111001", "00000011", "00001100", "00010101", "00011101", "00100101", "00101011", "00110001", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110000", "00101011", "00100100", "00011100", "00010100", "00001011", "00000010", "11111000", "11101111", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001010", "11001101", "11010011", "11011001", "11100000", "11101000", "11110001", "11111010", "00000011", "00001101", "00010101", "00011110", "00100101", "00101100", "00110001", "00110101", "00111000", "00111010", "00111001", "00111000", "00110100", "00110000", "00101010", "00100011", "00011100", "00010011", "00001010", "00000001", "11111000", "11101111", "11100110", "11011110", "11010111", "11010001", "11001100", "11001001", "11000111", "11000110", "11000111", "11001010", "11001110", "11010011", "11011001", "11100001", "11101001", "11110010", "11111011", "00000100", "00001101", "00010110", "00011110", "00100110", "00101100", "00110010", "00110110", "00111000", "00111010", "00111001", "00110111", "00110100", "00101111", "00101010", "00100011", "00011011", "00010010", "00001001", "00000000", "11110111", "11101110", "11100101", "11011101", "11010110", "11010001", "11001100", "11001001", "11000111", "11000110", "11001000", "11001010", "11001110", "11010100", "11011010", "11100010", "11101010", "11110011", "11111100", "00000101", "00001110", "00010111", "00011111", "00100111", "00101101", "00110010", "00110110", "00111001", "00111010", "00111001", "00110111", "00110100", "00101111", "00101001", "00100010", "00011010", "00010001", "00001000", "11111111", "11110110", "11101101", "11100100", "11011101", "11010110", "11010000", "11001100", "11001000", "11000111", "11000110", "11001000", "11001011", "11001111", "11010100", "11011011", "11100010", "11101011", "11110011", "11111101", "00000110", "00001111", "00011000", "00100000", "00100111", "00101101", "00110011", "00110110", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010001", "00001000", "11111110", "11110101", "11101100", "11100100", "11011100", "11010101", "11010000", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11001111", "11010101", "11011011", "11100011", "11101011", "11110100", "11111101", "00000111", "00010000", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010000", "00000111", "11111101", "11110100", "11101011", "11100011", "11011011", "11010101", "11001111", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11010000", "11010101", "11011100", "11100100", "11101100", "11110101", "11111110", "00001000", "00010001", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010", "00111001", "00110110", "00110011", "00101101", "00100111", "00100000", "00011000", "00001111", "00000110", "11111101", "11110011", "11101011", "11100010", "11011011", "11010100", "11001111", "11001011", "11001000", "11000110", "11000111", "11001000", "11001100", "11010000", "11010110", "11011101", "11100100", "11101101", "11110110", "11111111", "00001000", "00010001", "00011010", "00100010", "00101001", "00101111", "00110100", "00110111", "00111001", "00111010", "00111001", "00110110", "00110010", "00101101", "00100111", "00011111", "00010111", "00001110", "00000101", "11111100", "11110011", "11101010", "11100010", "11011010", "11010100", "11001110", "11001010", "11001000", "11000110", "11000111", "11001001", "11001100", "11010001", "11010110", "11011101", "11100101", "11101110", "11110111", "00000000", "00001001", "00010010", "00011011", "00100011", "00101010", "00101111", "00110100", "00110111", "00111001", "00111010", "00111000", "00110110", "00110010", "00101100", "00100110", "00011110", "00010110", "00001101", "00000100", "11111011", "11110010", "11101001", "11100001", "11011001", "11010011", "11001110", "11001010", "11000111", "11000110", "11000111", "11001001", "11001100", "11010001", "11010111", "11011110", "11100110", "11101111", "11111000", "00000001", "00001010", "00010011", "00011100", "00100011", "00101010", "00110000", "00110100", "00111000", "00111001", "00111010", "00111000", "00110101", "00110001", "00101100", "00100101", "00011110", "00010101", "00001101", "00000011", "11111010", "11110001", "11101000", "11100000", "11011001", "11010011", "11001101", "11001010", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11101111", "11111000", "00000010", "00001011", "00010100", "00011100", "00100100", "00101011", "00110000", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110001", "00101011", "00100101", "00011101", "00010101", "00001100", "00000011", "11111001", "11110000", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001001", "11001101", "11010010", "11011000", "11011111", "11100111", "11110000", "11111001", "00000011", "00001100", "00010101", "00011101", "00100101", "00101011", "00110001", "00110101", "00111000", "00111001", "00111001", "00111000", "00110101", "00110000", "00101011", "00100100", "00011100", "00010100", "00001011", "00000010", "11111000", "11101111", "11100111", "11011111", "11011000", "11010010", "11001101", "11001001", "11000111", "11000110", "11000111", "11001010", "11001101", "11010011", "11011001", "11100000", "11101000", "11110001", "11111010", "00000011", "00001101", "00010101", "00011110", "00100101", "00101100", "00110001", "00110101", "00111000", "00111010", "00111001", "00111000", "00110100", "00110000", "00101010", "00100011", "00011100", "00010011", "00001010", "00000001", "11111000", "11101111", "11100110", "11011110", "11010111", "11010001", "11001100", "11001001", "11000111", "11000110", "11000111", "11001010", "11001110", "11010011", "11011001", "11100001", "11101001", "11110010", "11111011", "00000100", "00001101", "00010110", "00011110", "00100110", "00101100", "00110010", "00110110", "00111000", "00111010", "00111001", "00110111", "00110100", "00101111", "00101010", "00100011", "00011011", "00010010", "00001001", "00000000", "11110111", "11101110", "11100101", "11011101", "11010110", "11010001", "11001100", "11001001", "11000111", "11000110", "11001000", "11001010", "11001110", "11010100", "11011010", "11100010", "11101010", "11110011", "11111100", "00000101", "00001110", "00010111", "00011111", "00100111", "00101101", "00110010", "00110110", "00111001", "00111010", "00111001", "00110111", "00110100", "00101111", "00101001", "00100010", "00011010", "00010001", "00001000", "11111111", "11110110", "11101101", "11100100", "11011101", "11010110", "11010000", "11001100", "11001000", "11000111", "11000110", "11001000", "11001011", "11001111", "11010100", "11011011", "11100010", "11101011", "11110011", "11111101", "00000110", "00001111", "00011000", "00100000", "00100111", "00101101", "00110011", "00110110", "00111001", "00111010", "00111001", "00110111", "00110011", "00101110", "00101000", "00100001", "00011001", "00010001", "00001000", "11111110", "11110101", "11101100", "11100100", "11011100", "11010101", "11010000", "11001011", "11001000", "11000111", "11000111", "11001000", "11001011", "11001111", "11010101", "11011011", "11100011", "11101011", "11110100", "11111101", "00000111", "00010000", "00011001", "00100001", "00101000", "00101110", "00110011", "00110111", "00111001", "00111010"));

end Inputs_test;

package body Inputs_Test is
end Inputs_Test;
