library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.ReSamplerTypes.all;

package outputs_test is

-- Declare constants

  constant outputs :outputarray := (
("00000000000000000000000000000000", "00000000000000000000000011110010", "11111111111111111111111001000111", "00000000000000000000000101001111", "11111111111111111111101100000101", "00000000000000000000000101011011", "11111111111111111111110001100010", "11111111111111111111111111001111", "00000000000000000000001001110010", "11111111111111111111001110011111", "00000000000000000000100011111001", "11111111111111111110101100111011", "00000000000000000000101110011100", "11111111111111111111010011000100", "11111111111111111111110111011101", "00000000000000000000111000010001", "11111111111111111101101100111000", "00000000000000000010101011000011", "11111111111111111100011011011101", "00000000000000000010111000000011", "11111111111111111110001100111111", "11111111111111111111100101101110", "00000000000000000011001100111001", "11111111111111111001101011100111", "00000000000000001000110011110111", "11111111111111110101111111110010", "00000000000000001001001101011010", "11111111111111111010101101100001", "11111111111111111110000011000000", "00000000000000001101101110011101", "11111111111111100001000100000011", "00000000000000111101011101110101", "11111111111101100111011110111110", "11111111111010100100001011000011", "11111111111111101111100000011001", "00000000000011110111010011000000", "00000000000111100010101010111111", "00000000001011011011001111000001", "00000000001110011010111111111001", "00000000010010000101110011110100", "00000000010100101010000011000100", "00000000010111010011001100100010", "00000000011001011001111010000011", "00000000011011001000001010001011", "00000000011100010101110001000010", "00000000011100101110001011000100", "00000000011101000100010101010101", "00000000011100001000010010101101", "00000000011010111001011010001111", "00000000011001101000000111000000", "00000000010111001001101110111100", "00000000010100100000001010101110", "00000000010001110101110101100000", "00000000001110100001101011100011", "00000000001011000100101011101100", "00000000000111000111010011011001", "00000000000011010000101110011001", "11111111111111100011010101110111", "11111111111011000111001000101111", "11111111110111100000010101011001", "11111111110011110111000111111100", "11111111110000001010100010000001", "11111111101101010000001010100000", "11111111101010001110101100111001", "11111111100111111101110110001011", "11111111100110001010100011111110", "11111111100100101110100100111100", "11111111100011100000010011000111", "11111111100011000001001010001100", "11111111100011100010000100100110", "11111111100011111010111101011011", "11111111100101011101010111000101", "11111111100111010011100001011110", "11111111101001001110000011100011", "11111111101100010010010111011000", "11111111101111001000000001100111", "11111111110010001110110100100000", "11111111110110000101110010111101", "11111111111001111101101011110111", "11111111111101110010110101001111", "00000000000001101010110010001110", "00000000000101011111110110110111", "00000000001001011000001100100110", "00000000001101001101000101100101", "00000000010000101000101001101010", "00000000010011101101101001000110", "00000000010110011000101101001111", "00000000011000110010011010100001", "00000000011010100101110110001111", "00000000011011101101010101111100", "00000000011100100001111110100010", "00000000011100111110111101110000", "00000000011100101111110000011100", "00000000011011101001101110000000", "00000000011010001001111000111010", "00000000011000001110100110000011", "00000000010110000010100110111110", "00000000010011011000101100101110", "00000000001111111101001010100100", "00000000001100100011011101000111", "00000000001000110110010111010011", "00000000000100111011100111100100", "00000000000001000110011011111001", "11111111111101010000000010101010", "11111111111001011001000010101101", "11111111110101100000100100011000", "11111111110010000011101111010101", "11111111101110100100010100100100", "11111111101011100010110011110010", "11111111101001001000000100101001", "11111111100110100011011100110010", "11111111100100111110111010111111", "11111111100100001001100110010101", "11111111100011001010100101010011", "11111111100011000111011000110111", "11111111100011111101101100001010", "11111111100100110011111110110111", "11111111100110010110001111111000", "11111111101000100001010000001000", "11111111101010100111100101001010", "11111111101101011010111001111100", "11111111110000110001011001011000", "11111111110100010111101110001110", "11111111111000010101001110010111", "11111111111100001000001000011111", "11111111111111111111110000111011", "00000000000011110111101001001110", "00000000000111101010100000101110", "00000000001011101000000000001101", "00000000001111001110010111110011", "00000000010010100100111001011000", "00000000010101011000010001000110", "00000000010111011110100111100011", "00000000011001101001100011100111", "00000000011011001011111111001011", "00000000011100000010010001100000", "00000000011100111000100110110001", "00000000011100110101011110000010", "00000000011011110110011110010000", "00000000011011000001001001000111", "00000000011001011100110001110110", "00000000010110111000000100011111", "00000000010100011101010101110000", "00000000010001011011111100111101", "00000000001101111100100001101101", "00000000001010011111101100011010", "00000000000110100111001100010010", "00000000000010110000001111010011", "11111111111110111001110011101101", "11111111111011000100101001010011", "11111111110111001001111011101000", "11111111110011011100110011000101", "11111111110000000011000011010010", "11111111101100100111100010110010", "11111111101001111101100010100110", "11111111100111110001100110011010", "11111111100101110110001110010001", "11111111100100010110011001000001", "11111111100011010000010011000100", "11111111100011000001000001001011", "11111111100011011101111010111000", "11111111100100010010100100111111", "11111111100101011010000010111111", "11111111100111001101011000111011", "11111111101001100111000111110000", "11111111101100010010001001011101", "11111111101111010111001000101000", "11111111110010110010101000011100", "11111111110110100111100000101000", "11111111111010011111111000010000", "11111111111110010100111100101110", "00000000000010001100110111011101", "00000000000110000010000011000110", "00000000001001111001110101110100", "00000000001101110000110111011001", "00000000010000110111110010001110", "00000000010011101101011010100010", "00000000010110110001101111010110", "00000000011000101100011000011111", "00000000011010100010011111000001", "00000000011100000100111010100000", "00000000011100011101111010000001", "00000000011100111110110001101100", "00000000011100011111101110110111", "00000000011011010001011101100111", "00000000011001110101100000101101", "00000000011000000010001001110101", "00000000010101110001011110111000", "00000000010010110000000001101011", "00000000001111110101011100100011", "00000000001100001001001010110111", "00000000001000011111010010110110", "00000000000100111001001100111001", "00000000000000011100011100010001", "11111111111100101111100100011111", "11111111111000111001000111101111", "11111111110100111010101110011110", "11111111110001011111011011000111", "11111111101110001000100110111011", "11111111101011100001010100110100", "11111111101000110101001011101111", "11111111100110011000011011101100", "11111111100101000111011000000010", "11111111100011110101100010110100", "11111111100010111111001010100001", "11111111100011001101001101011110", "11111111100011101110110001101111", "11111111100100110100010000010001", "11111111100110100111000001110100", "11111111101000101111001011011000", "11111111101011001111000100000000", "11111111101110000101001110110000", "11111111110001010110100110100001", "11111111110100110100001010011100", "11111111111000010000100000001100", "11111111111100001100011100111000", "00000000000000011111110000110110", "00000000000100011010000100001000", "00000000001000001111010001111010", "00000000001011111100011001010100", "00000000001111001110100000001010", "00000000010010101101101001101110", "00000000010101100101011011101011", "00000000010111101101100101101111", "00000000011001111011000010001001", "00000000011011100010001101110110", "00000000011100010110000010111000", "00000000011100100000100011101001", "00000000011100011111010111000110", "00000000011011111110001110011101", "00000000011010101100010100111101", "00000000011001001001110100101111", "00000000010110101111011111100010", "00000000010100001110001111010010", "00000000010001010111111101100101", "00000000001101110110011101000110", "00000000001010011011110100000100", "00000000000110100101111001010110", "00000000000010101111110100001100", "11111111111110100111001011011010", "11111111111010011011000111001010", "11111111110110101101011111101010", "11111111110010110100110001010101", "11111111101111011110001100110101", "11111111101100011110010000101000", "11111111101001101111101100011010", "11111111100111100011110000100000", "11111111100101011111110001001111", "11111111100100001001011010110100", "11111111100011011000101111111010", "11111111100011000000000000000001", "11111111100011011000101100110111", "11111111100100001001010111111011", "11111111100101011111101001001111", "11111111100111100011101000000100", "11111111101001101111100001001110", "11111111101100011110000001011010", "11111111101111011101111111101111", "11111111110010110100100000111010", "11111111110110101101001110100100", "11111111111010011010110110101101", "11111111111110100110110110010000", "00000000000010101111100010101100", "00000000000110100101100111100001", "00000000001010011011101000001000", "00000000001101110110001110100010", "00000000010001010111101011011110", "00000000010100001110000010110100", "00000000010110101111010011100110", "00000000011001001001101010010011", "00000000011010101100001101010100", "00000000011011111110001010000100", "00000000011100011111011000010100", "00000000011100100000100010000000", "00000000011100010110000111010111", "00000000011011100010010100110110", "00000000011001111011001011001110", "00000000010111101101101110111001", "00000000010101100101100101100111", "00000000010010101101111011000100", "00000000001111001110101110010101", "00000000001011111100100110010000", "00000000001000001111100010101011", "00000000000100011010010110100111", "00000000000000100000001000011001", "11111111111100001100101111000001", "11111111111000010000110001111110", "11111111110100110100011010000011", "11111111110001010110110101110011", "11111111101110000101011111011111", "11111111101011001111010001011011", "11111111101000101111010100110001", "11111111100110100111001100110101", "11111111100100110100011001010100", "11111111100011101110110101010001", "11111111100011001101010010010110", "11111111100010111111001011000000", "11111111100011110101011001111001", "11111111100101000111010100111100", "11111111100110011000010001100001", "11111111101000110100111010010110", "11111111101011100001001001110100", "11111111101110001000011011011000", "11111111110001011111001010011010", "11111111110100111010011100110110", "11111111111000111000110101011001", "11111111111100101111010110001010", "00000000000000011100001001000100", "00000000000100111000111101100111", "00000000001000011111000100010110", "00000000001100001000110111100100", "00000000001111110101001101001111", "00000000010010101111110101000100", "00000000010101110001010010011111", "00000000011000000010000000110001", "00000000011001110101011100000010", "00000000011011010001011011000100", "00000000011100011111101100111001", "00000000011100111110110101110100", "00000000011100011101111011011010", "00000000011100000101000010100101", "00000000011010100010101000111011", "00000000011000101100011110100010", "00000000010110110001111100011101", "00000000010011101101101000101000", "00000000010000110111111110011001", "00000000001101110001001011100000", "00000000001001111010001101000011", "00000000000110000010010100001001", "00000000000010001101001010110001", "11111111111110010101001101110010", "11111111111010100000001001001001", "11111111110110100111110011011010", "11111111110010110010111010011011", "11111111101111010111010110010110", "11111111101100010010010110111010", "11111111101001100111010010110001", "11111111100111001101100101011111", "11111111100101011010001001110001", "11111111100100010010101010000100", "11111111100011011110000001011110", "11111111100011000001000010010000", "11111111100011010000001111100100", "11111111100100010110010010000000", "11111111100101110110000111000110", "11111111100111110001011001111101", "11111111101001111101011001000010", "11111111101100100111010011010010", "11111111110000000010110101011100", "11111111110011011100100010111001", "11111111110111001001101000101101", "11111111111011000100011000011100", "11111111111110111001100100000111", "00000000000010101111111101010110", "00000000000110100110111101010011", "00000000001010011111011011101000", "00000000001101111100010000101011", "00000000010001011011101011011100", "00000000010100011101001100001110", "00000000010110110111111011010111", "00000000011001011100100011001110", "00000000011011000001000101000001", "00000000011011110110011001101011", "00000000011100110101011010101101", "00000000011100111000100111001001", "00000000011100000010010011110110", "00000000011011001100000001001001", "00000000011001101001110000001000", "00000000010111011110101111111000", "00000000010101011000011010110110", "00000000010010100101000110000100", "00000000001111001110100110101000", "00000000001011101000010001110010", "00000000000111101010110001101001", "00000000000011110111110111100001", "00000000000000000000001111000101", "11111111111100001000010110110010", "11111111111000010101011111010010", "11111111110100010111111111110011", "11111111110000110001101000001101", "11111111101101011011000110101000", "11111111101010100111101110111010", "11111111101000100001011000011101", "11111111100110010110011100011001", "11111111100100110100000000110101", "11111111100011111101101110100000", "11111111100011000111011001001111", "11111111100011001010100001111110", "11111111100100001001100001110000", "11111111100100111110110110111001", "11111111100110100011001110001010", "11111111101001000111111011100001", "11111111101011100010101010010000", "11111111101110100100000011000011", "11111111110010000011011110010011", "11111111110101100000010011100110", "11111111111001011000110011101110", "11111111111101001111110000101101", "00000000000001000110001100010011", "00000000000100111011010110101101", "00000000001000110110000100011000", "00000000001100100011001100111011", "00000000001111111100111100101110", "00000000010011011000011101001110", "00000000010110000010011101011010", "00000000011000001110011001100110", "00000000011010001001110001101111", "00000000011011101001100110111111", "00000000011100101111101100111100", "00000000011100111110111110110101", "00000000011100100010000101001000", "00000000011011101101011011000001", "00000000011010100101111101000001", "00000000011000110010100111000101", "00000000010110011000111000010000", "00000000010011101101110110100011", "00000000010000101000110111011000", "00000000001101001101010111100100", "00000000001001011000011111011000", "00000000000101100000000111110000", "00000000000001101011000011010010", "11111111111101110011001000100011", "11111111111001111101111100111010", "11111111110110000110001010001100", "11111111110010001111001000100111", "11111111101111001000001101110010", "11111111101100010010100101011110", "11111111101001001110010000101010", "11111111100111010011100111100001", "11111111100101011101100000111111", "11111111100011111011000101100000", "11111111100011100010000101111111", "11111111100011000001001110010100", "11111111100011100000010001001001", "11111111100100101110100010011001", "11111111100110001010011111010011", "11111111100111111101110110001011", "11111111101010001110100001001000", "11111111101101001111111110010101", "11111111110000001010100011011101", "11111111110011110110110101001001", "11111111110111100000101101001010", "11111111111011000110110011000111", "11111111111111100011100011101111", "00000000000011010000011011100001", "00000000000111000110111000010001", "00000000001011000101010001100010", "00000000001110100000100100111001", "00000000010001110111011001000101", "00000000010100011110101011001100", "00000000010111001010110100010001", "00000000011001100111100100010100", "00000000011010111000100111111110", "00000000011100001010011101001100", "00000000011101000000110101011111", "00000000011100110010110010100010", "00000000011100010001001110010001", "00000000011011001011101111101111", "00000000011001011000111110001100", "00000000010111010000110100101000", "00000000010100110000111100000000", "00000000010001111010110001010000", "00000000001110101001011001011111", "00000000001011001011110101100100", "00000000000111101111011111110100", "00000000000011110011100011001000", "11111111111111100000001111001010", "11111111111011100101111011111000", "11111111110111110000101110000110", "11111111110100000011100110101100", "11111111110000110001011111110110", "11111111101101010010010110010010", "11111111101010011010100100010101", "11111111101000010010011010010001", "11111111100110000100111101110111", "11111111100100011101110010001010", "11111111100011101001111101001000", "11111111100011011111011100010111", "11111111100011100000101000111010", "11111111100100000001110001100011", "11111111100101010011101011000011", "11111111100110110110001011010001", "11111111101001010000100000011110", "11111111101011110001110000101110", "11111111101110101000000010011011", "11111111110010001001100010111010", "11111111110101100100001011111100", "11111111111001011010000110101010", "11111111111101010000001011110100", "00000000000001011000110100100110", "00000000000101100100111000110110", "00000000001001010010100000010110", "00000000001101001011001110101011", "00000000010000100001110011001011", "00000000010011100001101111011000", "00000000010110010000010011100110", "00000000011000011100001111100000", "00000000011010100000001110110001", "00000000011011110110100101001100", "00000000011100100111010000000110", "00000000011100111111111111111111", "00000000011100100111010011001001", "00000000011011110110101000000101", "00000000011010100000010110110001", "00000000011000011100010111111100", "00000000010110010000011110110010", "00000000010011100001111110100110", "00000000010000100010000000010001", "00000000001101001011011111000110", "00000000001001010010110001011100", "00000000000101100101001001010011", "00000000000001011001001001110000", "11111111111101010000011101010100", "11111111111001011010011000011111", "11111111110101100100010111111000", "11111111110010001001110001011110", "11111111101110101000010100100010", "11111111101011110001111101001100", "11111111101001010000101100011010", "11111111100110110110010101101101", "11111111100101010011110010101100", "11111111100100000001110101111100", "11111111100011100000100111101100", "11111111100011011111011110000000", "11111111100011101001111000101001", "11111111100100011101101011001010", "11111111100110000100110100110010", "11111111101000010010010001000111", "11111111101010011010011010011001", "11111111101101010010000100111100", "11111111110000110001010001101011", "11111111110100000011011001110000", "11111111110111110000011101010101", "11111111111011100101101001011001", "11111111111111011111110111100111", "00000000000011110011010000111111", "00000000000111101111001110000010", "00000000001011001011100101111101", "00000000001110101001001010001101", "00000000010001111010100000100001", "00000000010100110000101110100101", "00000000010111010000101011001111", "00000000011001011000110011001011", "00000000011011001011100110101100", "00000000011100010001001010101111", "00000000011100110010101101101010", "00000000011101000000110101000000", "00000000011100001010100110000111", "00000000011010111000101011000100", "00000000011001100111101110011111", "00000000010111001011000101101010", "00000000010100011110110110001100", "00000000010001110111100100101000", "00000000001110100000110101100110", "00000000001011000101100011001010", "00000000000111000111001010100111", "00000000000011010000101001110110", "11111111111111100011110110111100", "11111111111011000111000010011001", "11111111110111100000111011101010", "11111111110011110111001000011100", "11111111110000001010110010110001", "11111111101101010000001010111100", "11111111101010001110101101100001", "11111111100111111101111111001111", "11111111100110001010100011111110", "11111111100100101110100100111100", "11111111100011100000010011000111", "11111111100011000001001010001100", "11111111100011100010000100100110", "11111111100011111010111101011011", "11111111100101011101010111000101", "11111111100111010011100001011110", "11111111101001001110000011100011", "11111111101100010010010111011000", "11111111101111001000000001100111", "11111111110010001110110100100000", "11111111110110000101110010111101", "11111111111001111101101011110111", "11111111111101110010110101001111", "00000000000001101010110010001110", "00000000000101011111110110110111", "00000000001001011000001100100110", "00000000001101001101000101100101", "00000000010000101000101001101010", "00000000010011101101101001000110", "00000000010110011000101101001111", "00000000011000110010011010100001", "00000000011010100101110110001111", "00000000011011101101010101111100", "00000000011100100001111110100010", "00000000011100111110111101110000", "00000000011100101111110000011100", "00000000011011101001101110000000", "00000000011010001001111000111010", "00000000011000001110100110000011", "00000000010110000010100110111110", "00000000010011011000101100101110", "00000000001111111101001010100100", "00000000001100100011011101000111", "00000000001000110110010111010011", "00000000000100111011100111100100", "00000000000001000110011011111001", "11111111111101010000000010101010", "11111111111001011001000010101101", "11111111110101100000100100011000", "11111111110010000011101111010101", "11111111101110100100010100100100", "11111111101011100010110011110010", "11111111101001001000000100101001", "11111111100110100011011100110010", "11111111100100111110111010111111", "11111111100100001001100110010101", "11111111100011001010100101010011", "11111111100011000111011000110111", "11111111100011111101101100001010", "11111111100100110011111110110111", "11111111100110010110001111111000", "11111111101000100001010000001000", "11111111101010100111100101001010", "11111111101101011010111001111100", "11111111110000110001011001011000", "11111111110100010111101110001110", "11111111111000010101001110010111", "11111111111100001000001000011111", "11111111111111111111110000111011", "00000000000011110111101001001110", "00000000000111101010100000101110", "00000000001011101000000000001101", "00000000001111001110010111110011", "00000000010010100100111001011000", "00000000010101011000010001000110", "00000000010111011110100111100011", "00000000011001101001100011100111", "00000000011011001011111111001011", "00000000011100000010010001100000", "00000000011100111000100110110001", "00000000011100110101011110000010", "00000000011011110110011110010000", "00000000011011000001001001000111", "00000000011001011100110001110110", "00000000010110111000000100011111", "00000000010100011101010101110000", "00000000010001011011111100111101", "00000000001101111100100001101101", "00000000001010011111101100011010", "00000000000110100111001100010010", "00000000000010110000001111010011", "11111111111110111001110011101101", "11111111111011000100101001010011", "11111111110111001001111011101000", "11111111110011011100110011000101", "11111111110000000011000011010010", "11111111101100100111100010110010", "11111111101001111101100010100110", "11111111100111110001100110011010", "11111111100101110110001110010001", "11111111100100010110011001000001", "11111111100011010000010011000100", "11111111100011000001000001001011", "11111111100011011101111010111000", "11111111100100010010100100111111", "11111111100101011010000010111111", "11111111100111001101011000111011", "11111111101001100111000111110000", "11111111101100010010001001011101", "11111111101111010111001000101000", "11111111110010110010101000011100", "11111111110110100111100000101000", "11111111111010011111111000010000", "11111111111110010100111100101110", "00000000000010001100110111011101", "00000000000110000010000011000110", "00000000001001111001110101110100", "00000000001101110000110111011001", "00000000010000110111110010001110", "00000000010011101101011010100010", "00000000010110110001101111010110", "00000000011000101100011000011111", "00000000011010100010011111000001", "00000000011100000100111010100000", "00000000011100011101111010000001", "00000000011100111110110001101100", "00000000011100011111101110110111", "00000000011011010001011101100111", "00000000011001110101100000101101", "00000000011000000010001001110101", "00000000010101110001011110111000", "00000000010010110000000001101011", "00000000001111110101011100100011", "00000000001100001001001010110111", "00000000001000011111010010110110", "00000000000100111001001100111001", "00000000000000011100011100010001", "11111111111100101111100100011111", "11111111111000111001000111101111", "11111111110100111010101110011110", "11111111110001011111011011000111", "11111111101110001000100110111011", "11111111101011100001010100110100", "11111111101000110101001011101111", "11111111100110011000011011101100", "11111111100101000111011000000010", "11111111100011110101100010110100", "11111111100010111111001010100001", "11111111100011001101001101011110", "11111111100011101110110001101111", "11111111100100110100010000010001", "11111111100110100111000001110100", "11111111101000101111001011011000", "11111111101011001111000100000000", "11111111101110000101001110110000", "11111111110001010110100110100001", "11111111110100110100001010011100", "11111111111000010000100000001100", "11111111111100001100011100111000", "00000000000000011111110000110110", "00000000000100011010000100001000", "00000000001000001111010001111010", "00000000001011111100011001010100", "00000000001111001110100000001010", "00000000010010101101101001101110", "00000000010101100101011011101011", "00000000010111101101100101101111", "00000000011001111011000010001001", "00000000011011100010001101110110", "00000000011100010110000010111000", "00000000011100100000100011101001", "00000000011100011111010111000110", "00000000011011111110001110011101", "00000000011010101100010100111101", "00000000011001001001110100101111", "00000000010110101111011111100010", "00000000010100001110001111010010", "00000000010001010111111101100101", "00000000001101110110011101000110", "00000000001010011011110100000100", "00000000000110100101111001010110", "00000000000010101111110100001100", "11111111111110100111001011011010", "11111111111010011011000111001010", "11111111110110101101011111101010", "11111111110010110100110001010101", "11111111101111011110001100110101", "11111111101100011110010000101000", "11111111101001101111101100011010", "11111111100111100011110000100000", "11111111100101011111110001001111", "11111111100100001001011010110100", "11111111100011011000101111111010", "11111111100011000000000000000001", "11111111100011011000101100110111", "11111111100100001001010111111011", "11111111100101011111101001001111", "11111111100111100011101000000100", "11111111101001101111100001001110", "11111111101100011110000001011010", "11111111101111011101111111101111", "11111111110010110100100000111010", "11111111110110101101001110100100", "11111111111010011010110110101101", "11111111111110100110110110010000", "00000000000010101111100010101100", "00000000000110100101100111100001", "00000000001010011011101000001000", "00000000001101110110001110100010", "00000000010001010111101011011110", "00000000010100001110000010110100", "00000000010110101111010011100110", "00000000011001001001101010010011", "00000000011010101100001101010100", "00000000011011111110001010000100", "00000000011100011111011000010100", "00000000011100100000100010000000", "00000000011100010110000111010111", "00000000011011100010010100110110", "00000000011001111011001011001110", "00000000010111101101101110111001", "00000000010101100101100101100111", "00000000010010101101111011000100", "00000000001111001110101110010101", "00000000001011111100100110010000", "00000000001000001111100010101011", "00000000000100011010010110100111", "00000000000000100000001000011001", "11111111111100001100101111000001", "11111111111000010000110001111110", "11111111110100110100011010000011", "11111111110001010110110101110011", "11111111101110000101011111011111", "11111111101011001111010001011011", "11111111101000101111010100110001", "11111111100110100111001100110101", "11111111100100110100011001010100", "11111111100011101110110101010001", "11111111100011001101010010010110", "11111111100010111111001011000000", "11111111100011110101011001111001", "11111111100101000111010100111100", "11111111100110011000010001100001", "11111111101000110100111010010110", "11111111101011100001001001110100", "11111111101110001000011011011000", "11111111110001011111001010011010", "11111111110100111010011100110110", "11111111111000111000110101011001", "11111111111100101111010110001010", "00000000000000011100001001000100", "00000000000100111000111101100111", "00000000001000011111000100010110", "00000000001100001000110111100100", "00000000001111110101001101001111", "00000000010010101111110101000100", "00000000010101110001010010011111", "00000000011000000010000000110001", "00000000011001110101011100000010", "00000000011011010001011011000100", "00000000011100011111101100111001", "00000000011100111110110101110100", "00000000011100011101111011011010", "00000000011100000101000010100101", "00000000011010100010101000111011", "00000000011000101100011110100010", "00000000010110110001111100011101", "00000000010011101101101000101000", "00000000010000110111111110011001", "00000000001101110001001011100000", "00000000001001111010001101000011", "00000000000110000010010100001001", "00000000000010001101001010110001", "11111111111110010101001101110010", "11111111111010100000001001001001", "11111111110110100111110011011010", "11111111110010110010111010011011", "11111111101111010111010110010110", "11111111101100010010010110111010", "11111111101001100111010010110001", "11111111100111001101100101011111", "11111111100101011010001001110001", "11111111100100010010101010000100", "11111111100011011110000001011110", "11111111100011000001000010010000", "11111111100011010000001111100100", "11111111100100010110010010000000", "11111111100101110110000111000110", "11111111100111110001011001111101", "11111111101001111101011001000010", "11111111101100100111010011010010", "11111111110000000010110101011100", "11111111110011011100100010111001", "11111111110111001001101000101101", "11111111111011000100011000011100", "11111111111110111001100100000111", "00000000000010101111111101010110", "00000000000110100110111101010011", "00000000001010011111011011101000", "00000000001101111100010000101011", "00000000010001011011101011011100", "00000000010100011101001100001110", "00000000010110110111111011010111", "00000000011001011100100011001110", "00000000011011000001000101000001", "00000000011011110110011001101011", "00000000011100110101011010101101", "00000000011100111000100111001001", "00000000011100000010010011110110", "00000000011011001100000001001001", "00000000011001101001110000001000", "00000000010111011110101111111000", "00000000010101011000011010110110", "00000000010010100101000110000100", "00000000001111001110100110101000", "00000000001011101000010001110010", "00000000000111101010110001101001", "00000000000011110111110111100001", "00000000000000000000001111000101", "11111111111100001000010110110010", "11111111111000010101011111010010", "11111111110100010111111111110011", "11111111110000110001101000001101", "11111111101101011011000110101000", "11111111101010100111101110111010", "11111111101000100001011000011101", "11111111100110010110011100011001", "11111111100100110100000000110101", "11111111100011111101101110100000", "11111111100011000111011001001111", "11111111100011001010100001111110", "11111111100100001001100001110000", "11111111100100111110110110111001", "11111111100110100011001110001010", "11111111101001000111111011100001", "11111111101011100010101010010000", "11111111101110100100000011000011", "11111111110010000011011110010011", "11111111110101100000010011100110", "11111111111001011000110011101110", "11111111111101001111110000101101", "00000000000001000110001100010011", "00000000000100111011010110101101", "00000000001000110110000100011000", "00000000001100100011001100111011", "00000000001111111100111100101110", "00000000010011011000011101001110", "00000000010110000010011101011010", "00000000011000001110011001100110", "00000000011010001001110001101111", "00000000011011101001100110111111", "00000000011100101111101100111100", "00000000011100111110111110110101", "00000000011100100010000101001000", "00000000011011101101011011000001", "00000000011010100101111101000001", "00000000011000110010100111000101", "00000000010110011000111000010000", "00000000010011101101110110100011", "00000000010000101000110111011000", "00000000001101001101010111100100", "00000000001001011000011111011000", "00000000000101100000000111110000", "00000000000001101011000011010010", "11111111111101110011001000100011", "11111111111001111101111100111010", "11111111110110000110001010001100", "11111111110010001111001000100111", "11111111101111001000001101110010", "11111111101100010010100101011110", "11111111101001001110010000101010", "11111111100111010011100111100001", "11111111100101011101100000111111", "11111111100011111011000101100000", "11111111100011100010000101111111", "11111111100011000001001110010100", "11111111100011100000010001001001", "11111111100100101110100010011001", "11111111100110001010011111010011", "11111111100111111101110110001011", "11111111101010001110100001001000", "11111111101101001111111110010101", "11111111110000001010100011011101", "11111111110011110110110101001001", "11111111110111100000101101001010", "11111111111011000110110011000111", "11111111111111100011100011101111", "00000000000011010000011011100001", "00000000000111000110111000010001", "00000000001011000101010001100010", "00000000001110100000100100111001", "00000000010001110111011001000101", "00000000010100011110101011001100", "00000000010111001010110100010001", "00000000011001100111100100010100", "00000000011010111000100111111110", "00000000011100001010011101001100", "00000000011101000000110101011111", "00000000011100110010110010100010", "00000000011100010001001110010001", "00000000011011001011101111101111", "00000000011001011000111110001100", "00000000010111010000110100101000", "00000000010100110000111100000000", "00000000010001111010110001010000", "00000000001110101001011001011111", "00000000001011001011110101100100", "00000000000111101111011111110100", "00000000000011110011100011001000", "11111111111111100000001111001010", "11111111111011100101111011111000", "11111111110111110000101110000110", "11111111110100000011100110101100", "11111111110000110001011111110110", "11111111101101010010010110010010", "11111111101010011010100100010101", "11111111101000010010011010010001", "11111111100110000100111101110111", "11111111100100011101110010001010", "11111111100011101001111101001000", "11111111100011011111011100010111", "11111111100011100000101000111010", "11111111100100000001110001100011", "11111111100101010011101011000011", "11111111100110110110001011010001", "11111111101001010000100000011110", "11111111101011110001110000101110", "11111111101110101000000010011011", "11111111110010001001100010111010", "11111111110101100100001011111100", "11111111111001011010000110101010", "11111111111101010000001011110100", "00000000000001011000110100100110", "00000000000101100100111000110110", "00000000001001010010100000010110", "00000000001101001011001110101011", "00000000010000100001110011001011", "00000000010011100001101111011000", "00000000010110010000010011100110", "00000000011000011100001111100000", "00000000011010100000001110110001", "00000000011011110110100101001100", "00000000011100100111010000000110", "00000000011100111111111111111111", "00000000011100100111010011001001", "00000000011011110110101000000101", "00000000011010100000010110110001", "00000000011000011100010111111100", "00000000010110010000011110110010", "00000000010011100001111110100110", "00000000010000100010000000010001", "00000000001101001011011111000110", "00000000001001010010110001011100", "00000000000101100101001001010011", "00000000000001011001001001110000", "11111111111101010000011101010100", "11111111111001011010011000011111", "11111111110101100100010111111000", "11111111110010001001110001011110", "11111111101110101000010100100010", "11111111101011110001111101001100", "11111111101001010000101100011010", "11111111100110110110010101101101", "11111111100101010011110010101100", "11111111100100000001110101111100", "11111111100011100000100111101100", "11111111100011011111011110000000", "11111111100011101001111000101001", "11111111100100011101101011001010", "11111111100110000100110100110010", "11111111101000010010010001000111", "11111111101010011010011010011001", "11111111101101010010000100111100", "11111111110000110001010001101011", "11111111110100000011011001110000", "11111111110111110000011101010101", "11111111111011100101101001011001", "11111111111111011111110111100111", "00000000000011110011010000111111", "00000000000111101111001110000010", "00000000001011001011100101111101", "00000000001110101001001010001101", "00000000010001111010100000100001", "00000000010100110000101110100101", "00000000010111010000101011001111", "00000000011001011000110011001011", "00000000011011001011100110101100", "00000000011100010001001010101111", "00000000011100110010101101101010", "00000000011101000000110101000000", "00000000011100001010100110000111", "00000000011010111000101011000100", "00000000011001100111101110011111", "00000000010111001011000101101010", "00000000010100011110110110001100", "00000000010001110111100100101000", "00000000001110100000110101100110", "00000000001011000101100011001010", "00000000000111000111001010100111", "00000000000011010000101001110110", "11111111111111100011110110111100", "11111111111011000111000010011001", "11111111110111100000111011101010", "11111111110011110111001000011100", "11111111110000001010110010110001", "11111111101101010000001010111100", "11111111101010001110101101100001", "11111111100111111101111111001111", "11111111100110001010100011111110", "11111111100100101110100100111100", "11111111100011100000010011000111", "11111111100011000001001010001100", "11111111100011100010000100100110", "11111111100011111010111101011011", "11111111100101011101010111000101", "11111111100111010011100001011110", "11111111101001001110000011100011", "11111111101100010010010111011000", "11111111101111001000000001100111", "11111111110010001110110100100000", "11111111110110000101110010111101", "11111111111001111101101011110111", "11111111111101110010110101001111", "00000000000001101010110010001110", "00000000000101011111110110110111", "00000000001001011000001100100110", "00000000001101001101000101100101", "00000000010000101000101001101010", "00000000010011101101101001000110", "00000000010110011000101101001111", "00000000011000110010011010100001", "00000000011010100101110110001111", "00000000011011101101010101111100", "00000000011100100001111110100010", "00000000011100111110111101110000", "00000000011100101111110000011100", "00000000011011101001101110000000", "00000000011010001001111000111010", "00000000011000001110100110000011", "00000000010110000010100110111110", "00000000010011011000101100101110", "00000000001111111101001010100100", "00000000001100100011011101000111", "00000000001000110110010111010011", "00000000000100111011100111100100", "00000000000001000110011011111001", "11111111111101010000000010101010", "11111111111001011001000010101101", "11111111110101100000100100011000", "11111111110010000011101111010101", "11111111101110100100010100100100", "11111111101011100010110011110010", "11111111101001001000000100101001", "11111111100110100011011100110010", "11111111100100111110111010111111", "11111111100100001001100110010101", "11111111100011001010100101010011", "11111111100011000111011000110111", "11111111100011111101101100001010", "11111111100100110011111110110111", "11111111100110010110001111111000", "11111111101000100001010000001000", "11111111101010100111100101001010", "11111111101101011010111001111100", "11111111110000110001011001011000", "11111111110100010111101110001110", "11111111111000010101001110010111", "11111111111100001000001000011111", "11111111111111111111110000111011", "00000000000011110111101001001110", "00000000000111101010100000101110", "00000000001011101000000000001101", "00000000001111001110010111110011", "00000000010010100100111001011000", "00000000010101011000010001000110", "00000000010111011110100111100011", "00000000011001101001100011100111", "00000000011011001011111111001011", "00000000011100000010010001100000", "00000000011100111000100110110001", "00000000011100110101011110000010", "00000000011011110110011110010000", "00000000011011000001001001000111", "00000000011001011100110001110110", "00000000010110111000000100011111", "00000000010100011101010101110000", "00000000010001011011111100111101", "00000000001101111100100001101101", "00000000001010011111101100011010", "00000000000110100111001100010010", "00000000000010110000001111010011", "11111111111110111001110011101101", "11111111111011000100101001010011", "11111111110111001001111011101000", "11111111110011011100110011000101", "11111111110000000011000011010010", "11111111101100100111100010110010", "11111111101001111101100010100110", "11111111100111110001100110011010", "11111111100101110110001110010001", "11111111100100010110011001000001", "11111111100011010000010011000100", "11111111100011000001000001001011", "11111111100011011101111010111000", "11111111100100010010100100111111", "11111111100101011010000010111111", "11111111100111001101011000111011", "11111111101001100111000111110000", "11111111101100010010001001011101", "11111111101111010111001000101000", "11111111110010110010101000011100", "11111111110110100111100000101000", "11111111111010011111111000010000", "11111111111110010100111100101110", "00000000000010001100110111011101", "00000000000110000010000011000110", "00000000001001111001110101110100", "00000000001101110000110111011001", "00000000010000110111110010001110", "00000000010011101101011010100010", "00000000010110110001101111010110", "00000000011000101100011000011111", "00000000011010100010011111000001", "00000000011100000100111010100000", "00000000011100011101111010000001", "00000000011100111110110001101100", "00000000011100011111101110110111", "00000000011011010001011101100111", "00000000011001110101100000101101", "00000000011000000010001001110101", "00000000010101110001011110111000", "00000000010010110000000001101011", "00000000001111110101011100100011", "00000000001100001001001010110111", "00000000001000011111010010110110", "00000000000100111001001100111001", "00000000000000011100011100010001", "11111111111100101111100100011111", "11111111111000111001000111101111", "11111111110100111010101110011110", "11111111110001011111011011000111", "11111111101110001000100110111011", "11111111101011100001010100110100", "11111111101000110101001011101111", "11111111100110011000011011101100", "11111111100101000111011000000010", "11111111100011110101100010110100", "11111111100010111111001010100001", "11111111100011001101001101011110", "11111111100011101110110001101111", "11111111100100110100010000010001", "11111111100110100111000001110100", "11111111101000101111001011011000", "11111111101011001111000100000000", "11111111101110000101001110110000", "11111111110001010110100110100001", "11111111110100110100001010011100", "11111111111000010000100000001100", "11111111111100001100011100111000", "00000000000000011111110000110110", "00000000000100011010000100001000", "00000000001000001111010001111010", "00000000001011111100011001010100", "00000000001111001110100000001010", "00000000010010101101101001101110", "00000000010101100101011011101011", "00000000010111101101100101101111", "00000000011001111011000010001001", "00000000011011100010001101110110", "00000000011100010110000010111000", "00000000011100100000100011101001", "00000000011100011111010111000110", "00000000011011111110001110011101", "00000000011010101100010100111101", "00000000011001001001110100101111", "00000000010110101111011111100010", "00000000010100001110001111010010", "00000000010001010111111101100101", "00000000001101110110011101000110", "00000000001010011011110100000100", "00000000000110100101111001010110", "00000000000010101111110100001100", "11111111111110100111001011011010", "11111111111010011011000111001010", "11111111110110101101011111101010", "11111111110010110100110001010101", "11111111101111011110001100110101", "11111111101100011110010000101000", "11111111101001101111101100011010", "11111111100111100011110000100000", "11111111100101011111110001001111", "11111111100100001001011010110100", "11111111100011011000101111111010", "11111111100011000000000000000001", "11111111100011011000101100110111", "11111111100100001001010111111011", "11111111100101011111101001001111", "11111111100111100011101000000100", "11111111101001101111100001001110", "11111111101100011110000001011010", "11111111101111011101111111101111", "11111111110010110100100000111010", "11111111110110101101001110100100", "11111111111010011010110110101101", "11111111111110100110110110010000", "00000000000010101111100010101100", "00000000000110100101100111100001", "00000000001010011011101000001000", "00000000001101110110001110100010", "00000000010001010111101011011110", "00000000010100001110000010110100", "00000000010110101111010011100110", "00000000011001001001101010010011", "00000000011010101100001101010100", "00000000011011111110001010000100", "00000000011100011111011000010100", "00000000011100100000100010000000", "00000000011100010110000111010111", "00000000011011100010010100110110", "00000000011001111011001011001110", "00000000010111101101101110111001", "00000000010101100101100101100111", "00000000010010101101111011000100", "00000000001111001110101110010101", "00000000001011111100100110010000", "00000000001000001111100010101011", "00000000000100011010010110100111", "00000000000000100000001000011001", "11111111111100001100101111000001", "11111111111000010000110001111110", "11111111110100110100011010000011", "11111111110001010110110101110011", "11111111101110000101011111011111", "11111111101011001111010001011011", "11111111101000101111010100110001", "11111111100110100111001100110101", "11111111100100110100011001010100", "11111111100011101110110101010001", "11111111100011001101010010010110", "11111111100010111111001011000000", "11111111100011110101011001111001", "11111111100101000111010100111100", "11111111100110011000010001100001", "11111111101000110100111010010110", "11111111101011100001001001110100", "11111111101110001000011011011000", "11111111110001011111001010011010", "11111111110100111010011100110110", "11111111111000111000110101011001", "11111111111100101111010110001010", "00000000000000011100001001000100", "00000000000100111000111101100111", "00000000001000011111000100010110", "00000000001100001000110111100100", "00000000001111110101001101001111", "00000000010010101111110101000100", "00000000010101110001010010011111", "00000000011000000010000000110001", "00000000011001110101011100000010", "00000000011011010001011011000100", "00000000011100011111101100111001", "00000000011100111110110101110100", "00000000011100011101111011011010", "00000000011100000101000010100101", "00000000011010100010101000111011", "00000000011000101100011110100010", "00000000010110110001111100011101", "00000000010011101101101000101000", "00000000010000110111111110011001", "00000000001101110001001011100000", "00000000001001111010001101000011", "00000000000110000010010100001001", "00000000000010001101001010110001", "11111111111110010101001101110010", "11111111111010100000001001001001", "11111111110110100111110011011010", "11111111110010110010111010011011", "11111111101111010111010110010110", "11111111101100010010010110111010", "11111111101001100111010010110001", "11111111100111001101100101011111", "11111111100101011010001001110001", "11111111100100010010101010000100", "11111111100011011110000001011110", "11111111100011000001000010010000", "11111111100011010000001111100100", "11111111100100010110010010000000", "11111111100101110110000111000110", "11111111100111110001011001111101", "11111111101001111101011001000010", "11111111101100100111010011010010", "11111111110000000010110101011100", "11111111110011011100100010111001", "11111111110111001001101000101101", "11111111111011000100011000011100", "11111111111110111001100100000111", "00000000000010101111111101010110", "00000000000110100110111101010011", "00000000001010011111011011101000", "00000000001101111100010000101011", "00000000010001011011101011011100", "00000000010100011101001100001110", "00000000010110110111111011010111", "00000000011001011100100011001110", "00000000011011000001000101000001", "00000000011011110110011001101011", "00000000011100110101011010101101", "00000000011100111000100111001001", "00000000011100000010010011110110", "00000000011011001100000001001001", "00000000011001101001110000001000", "00000000010111011110101111111000", "00000000010101011000011010110110", "00000000010010100101000110000100", "00000000001111001110100110101000", "00000000001011101000010001110010", "00000000000111101010110001101001", "00000000000011110111110111100001", "00000000000000000000001111000101", "11111111111100001000010110110010", "11111111111000010101011111010010", "11111111110100010111111111110011", "11111111110000110001101000001101", "11111111101101011011000110101000", "11111111101010100111101110111010", "11111111101000100001011000011101", "11111111100110010110011100011001", "11111111100100110100000000110101", "11111111100011111101101110100000", "11111111100011000111011001001111", "11111111100011001010100001111110", "11111111100100001001100001110000", "11111111100100111110110110111001", "11111111100110100011001110001010", "11111111101001000111111011100001", "11111111101011100010101010010000", "11111111101110100100000011000011", "11111111110010000011011110010011", "11111111110101100000010011100110", "11111111111001011000110011101110", "11111111111101001111110000101101", "00000000000001000110001100010011", "00000000000100111011010110101101", "00000000001000110110000100011000", "00000000001100100011001100111011", "00000000001111111100111100101110", "00000000010011011000011101001110", "00000000010110000010011101011010", "00000000011000001110011001100110", "00000000011010001001110001101111", "00000000011011101001100110111111", "00000000011100101111101100111100", "00000000011100111110111110110101", "00000000011100100010000101001000", "00000000011011101101011011000001", "00000000011010100101111101000001", "00000000011000110010100111000101", "00000000010110011000111000010000", "00000000010011101101110110100011", "00000000010000101000110111011000", "00000000001101001101010111100100", "00000000001001011000011111011000", "00000000000101100000000111110000", "00000000000001101011000011010010", "11111111111101110011001000100011", "11111111111001111101111100111010", "11111111110110000110001010001100", "11111111110010001111001000100111", "11111111101111001000001101110010", "11111111101100010010100101011110", "11111111101001001110010000101010", "11111111100111010011100111100001", "11111111100101011101100000111111", "11111111100011111011000101100000", "11111111100011100010000101111111", "11111111100011000001001110010100", "11111111100011100000010001001001", "11111111100100101110100010011001", "11111111100110001010011111010011", "11111111100111111101110110001011", "11111111101010001110100001001000", "11111111101101001111111110010101", "11111111110000001010100011011101", "11111111110011110110110101001001", "11111111110111100000101101001010", "11111111111011000110110011000111", "11111111111111100011100011101111", "00000000000011010000011011100001", "00000000000111000110111000010001", "00000000001011000101010001100010", "00000000001110100000100100111001", "00000000010001110111011001000101", "00000000010100011110101011001100", "00000000010111001010110100010001", "00000000011001100111100100010100", "00000000011010111000100111111110", "00000000011100001010011101001100", "00000000011101000000110101011111", "00000000011100110010110010100010", "00000000011100010001001110010001", "00000000011011001011101111101111", "00000000011001011000111110001100", "00000000010111010000110100101000", "00000000010100110000111100000000", "00000000010001111010110001010000", "00000000001110101001011001011111", "00000000001011001011110101100100", "00000000000111101111011111110100", "00000000000011110011100011001000", "11111111111111100000001111001010", "11111111111011100101111011111000", "11111111110111110000101110000110", "11111111110100000011100110101100", "11111111110000110001011111110110", "11111111101101010010010110010010", "11111111101010011010100100010101", "11111111101000010010011010010001", "11111111100110000100111101110111", "11111111100100011101110010001010", "11111111100011101001111101001000", "11111111100011011111011100010111", "11111111100011100000101000111010", "11111111100100000001110001100011", "11111111100101010011101011000011", "11111111100110110110001011010001", "11111111101001010000100000011110", "11111111101011110001110000101110", "11111111101110101000000010011011", "11111111110010001001100010111010", "11111111110101100100001011111100", "11111111111001011010000110101010", "11111111111101010000001011110100", "00000000000001011000110100100110", "00000000000101100100111000110110", "00000000001001010010100000010110", "00000000001101001011001110101011", "00000000010000100001110011001011", "00000000010011100001101111011000", "00000000010110010000010011100110", "00000000011000011100001111100000", "00000000011010100000001110110001", "00000000011011110110100101001100", "00000000011100100111010000000110", "00000000011100111111111111111111", "00000000011100100111010011001001", "00000000011011110110101000000101", "00000000011010100000010110110001", "00000000011000011100010111111100", "00000000010110010000011110110010", "00000000010011100001111110100110", "00000000010000100010000000010001", "00000000001101001011011111000110", "00000000001001010010110001011100", "00000000000101100101001001010011", "00000000000001011001001001110000", "11111111111101010000011101010100", "11111111111001011010011000011111", "11111111110101100100010111111000", "11111111110010001001110001011110", "11111111101110101000010100100010", "11111111101011110001111101001100", "11111111101001010000101100011010", "11111111100110110110010101101101", "11111111100101010011110010101100", "11111111100100000001110101111100", "11111111100011100000100111101100", "11111111100011011111011110000000", "11111111100011101001111000101001", "11111111100100011101101011001010", "11111111100110000100110100110010", "11111111101000010010010001000111", "11111111101010011010011010011001", "11111111101101010010000100111100", "11111111110000110001010001101011", "11111111110100000011011001110000", "11111111110111110000011101010101", "11111111111011100101101001011001", "11111111111111011111110111100111", "00000000000011110011010000111111", "00000000000111101111001110000010", "00000000001011001011100101111101", "00000000001110101001001010001101", "00000000010001111010100000100001", "00000000010100110000101110100101", "00000000010111010000101011001111", "00000000011001011000110011001011", "00000000011011001011100110101100", "00000000011100010001001010101111", "00000000011100110010101101101010", "00000000011101000000110101000000", "00000000011100001010100110000111", "00000000011010111000101011000100", "00000000011001100111101110011111", "00000000010111001011000101101010", "00000000010100011110110110001100", "00000000010001110111100100101000", "00000000001110100000110101100110", "00000000001011000101100011001010", "00000000000111000111001010100111", "00000000000011010000101001110110", "11111111111111100011110110111100", "11111111111011000111000010011001", "11111111110111100000111011101010", "11111111110011110111001000011100", "11111111110000001010110010110001", "11111111101101010000001010111100", "11111111101010001110101101100001", "11111111100111111101111111001111", "11111111100110001010100011111110", "11111111100100101110100100111100", "11111111100011100000010011000111", "11111111100011000001001010001100", "11111111100011100010000100100110", "11111111100011111010111101011011", "11111111100101011101010111000101", "11111111100111010011100001011110", "11111111101001001110000011100011", "11111111101100010010010111011000", "11111111101111001000000001100111", "11111111110010001110110100100000", "11111111110110000101110010111101", "11111111111001111101101011110111", "11111111111101110010110101001111", "00000000000001101010110010001110", "00000000000101011111110110110111", "00000000001001011000001100100110", "00000000001101001101000101100101", "00000000010000101000101001101010", "00000000010011101101101001000110", "00000000010110011000101101001111", "00000000011000110010011010100001", "00000000011010100101110110001111", "00000000011011101101010101111100", "00000000011100100001111110100010", "00000000011100111110111101110000", "00000000011100101111110000011100", "00000000011011101001101110000000", "00000000011010001001111000111010", "00000000011000001110100110000011", "00000000010110000010100110111110", "00000000010011011000101100101110", "00000000001111111101001010100100", "00000000001100100011011101000111", "00000000001000110110010111010011", "00000000000100111011100111100100", "00000000000001000110011011111001", "11111111111101010000000010101010", "11111111111001011001000010101101", "11111111110101100000100100011000", "11111111110010000011101111010101", "11111111101110100100010100100100", "11111111101011100010110011110010", "11111111101001001000000100101001", "11111111100110100011011100110010", "11111111100100111110111010111111", "11111111100100001001100110010101", "11111111100011001010100101010011", "11111111100011000111011000110111", "11111111100011111101101100001010", "11111111100100110011111110110111", "11111111100110010110001111111000", "11111111101000100001010000001000", "11111111101010100111100101001010", "11111111101101011010111001111100", "11111111110000110001011001011000", "11111111110100010111101110001110", "11111111111000010101001110010111", "11111111111100001000001000011111", "11111111111111111111110000111011", "00000000000011110111101001001110", "00000000000111101010100000101110", "00000000001011101000000000001101", "00000000001111001110010111110011", "00000000010010100100111001011000", "00000000010101011000010001000110", "00000000010111011110100111100011", "00000000011001101001100011100111", "00000000011011001011111111001011", "00000000011100000010010001100000", "00000000011100111000100110110001", "00000000011100110101011110000010", "00000000011011110110011110010000", "00000000011011000001001001000111", "00000000011001011100110001110110", "00000000010110111000000100011111", "00000000010100011101010101110000", "00000000010001011011111100111101", "00000000001101111100100001101101", "00000000001010011111101100011010", "00000000000110100111001100010010", "00000000000010110000001111010011", "11111111111110111001110011101101", "11111111111011000100101001010011", "11111111110111001001111011101000", "11111111110011011100110011000101", "11111111110000000011000011010010", "11111111101100100111100010110010", "11111111101001111101100010100110", "11111111100111110001100110011010", "11111111100101110110001110010001", "11111111100100010110011001000001", "11111111100011010000010011000100", "11111111100011000001000001001011", "11111111100011011101111010111000", "11111111100100010010100100111111", "11111111100101011010000010111111", "11111111100111001101011000111011", "11111111101001100111000111110000", "11111111101100010010001001011101", "11111111101111010111001000101000", "11111111110010110010101000011100", "11111111110110100111100000101000", "11111111111010011111111000010000", "11111111111110010100111100101110", "00000000000010001100110111011101", "00000000000110000010000011000110", "00000000001001111001110101110100", "00000000001101110000110111011001", "00000000010000110111110010001110", "00000000010011101101011010100010", "00000000010110110001101111010110", "00000000011000101100011000011111", "00000000011010100010011111000001", "00000000011100000100111010100000", "00000000011100011101111010000001", "00000000011100111110110001101100", "00000000011100011111101110110111", "00000000011011010001011101100111", "00000000011001110101100000101101", "00000000011000000010001001110101", "00000000010101110001011110111000", "00000000010010110000000001101011", "00000000001111110101011100100011", "00000000001100001001001010110111", "00000000001000011111010010110110", "00000000000100111001001100111001", "00000000000000011100011100010001", "11111111111100101111100100011111", "11111111111000111001000111101111", "11111111110100111010101110011110", "11111111110001011111011011000111", "11111111101110001000100110111011", "11111111101011100001010100110100", "11111111101000110101001011101111", "11111111100110011000011011101100", "11111111100101000111011000000010", "11111111100011110101100010110100", "11111111100010111111001010100001", "11111111100011001101001101011110", "11111111100011101110110001101111", "11111111100100110100010000010001", "11111111100110100111000001110100", "11111111101000101111001011011000", "11111111101011001111000100000000", "11111111101110000101001110110000", "11111111110001010110100110100001", "11111111110100110100001010011100", "11111111111000010000100000001100", "11111111111100001100011100111000", "00000000000000011111110000110110", "00000000000100011010000100001000", "00000000001000001111010001111010", "00000000001011111100011001010100", "00000000001111001110100000001010", "00000000010010101101101001101110", "00000000010101100101011011101011", "00000000010111101101100101101111", "00000000011001111011000010001001", "00000000011011100010001101110110", "00000000011100010110000010111000", "00000000011100100000100011101001", "00000000011100011111010111000110", "00000000011011111110001110011101", "00000000011010101100010100111101", "00000000011001001001110100101111", "00000000010110101111011111100010", "00000000010100001110001111010010", "00000000010001010111111101100101", "00000000001101110110011101000110", "00000000001010011011110100000100", "00000000000110100101111001010110", "00000000000010101111110100001100", "11111111111110100111001011011010", "11111111111010011011000111001010", "11111111110110101101011111101010", "11111111110010110100110001010101", "11111111101111011110001100110101", "11111111101100011110010000101000", "11111111101001101111101100011010", "11111111100111100011110000100000", "11111111100101011111110001001111", "11111111100100001001011010110100", "11111111100011011000101111111010", "11111111100011000000000000000001", "11111111100011011000101100110111", "11111111100100001001010111111011", "11111111100101011111101001001111", "11111111100111100011101000000100", "11111111101001101111100001001110", "11111111101100011110000001011010", "11111111101111011101111111101111", "11111111110010110100100000111010", "11111111110110101101001110100100", "11111111111010011010110110101101", "11111111111110100110110110010000", "00000000000010101111100010101100", "00000000000110100101100111100001", "00000000001010011011101000001000", "00000000001101110110001110100010", "00000000010001010111101011011110", "00000000010100001110000010110100", "00000000010110101111010011100110", "00000000011001001001101010010011", "00000000011010101100001101010100", "00000000011011111110001010000100", "00000000011100011111011000010100", "00000000011100100000100010000000", "00000000011100010110000111010111", "00000000011011100010010100110110", "00000000011001111011001011001110", "00000000010111101101101110111001", "00000000010101100101100101100111", "00000000010010101101111011000100", "00000000001111001110101110010101", "00000000001011111100100110010000", "00000000001000001111100010101011", "00000000000100011010010110100111", "00000000000000100000001000011001", "11111111111100001100101111000001", "11111111111000010000110001111110", "11111111110100110100011010000011", "11111111110001010110110101110011", "11111111101110000101011111011111", "11111111101011001111010001011011", "11111111101000101111010100110001", "11111111100110100111001100110101", "11111111100100110100011001010100", "11111111100011101110110101010001", "11111111100011001101010010010110", "11111111100010111111001011000000", "11111111100011110101011001111001", "11111111100101000111010100111100", "11111111100110011000010001100001", "11111111101000110100111010010110", "11111111101011100001001001110100", "11111111101110001000011011011000", "11111111110001011111001010011010", "11111111110100111010011100110110", "11111111111000111000110101011001", "11111111111100101111010110001010", "00000000000000011100001001000100", "00000000000100111000111101100111", "00000000001000011111000100010110", "00000000001100001000110111100100", "00000000001111110101001101001111", "00000000010010101111110101000100", "00000000010101110001010010011111", "00000000011000000010000000110001", "00000000011001110101011100000010", "00000000011011010001011011000100", "00000000011100011111101100111001", "00000000011100111110110101110100", "00000000011100011101111011011010", "00000000011100000101000010100101", "00000000011010100010101000111011", "00000000011000101100011110100010", "00000000010110110001111100011101", "00000000010011101101101000101000", "00000000010000110111111110011001", "00000000001101110001001011100000", "00000000001001111010001101000011", "00000000000110000010010100001001", "00000000000010001101001010110001", "11111111111110010101001101110010", "11111111111010100000001001001001", "11111111110110100111110011011010", "11111111110010110010111010011011", "11111111101111010111010110010110", "11111111101100010010010110111010", "11111111101001100111010010110001", "11111111100111001101100101011111", "11111111100101011010001001110001", "11111111100100010010101010000100", "11111111100011011110000001011110", "11111111100011000001000010010000", "11111111100011010000001111100100", "11111111100100010110010010000000", "11111111100101110110000111000110", "11111111100111110001011001111101", "11111111101001111101011001000010", "11111111101100100111010011010010", "11111111110000000010110101011100", "11111111110011011100100010111001", "11111111110111001001101000101101", "11111111111011000100011000011100", "11111111111110111001100100000111", "00000000000010101111111101010110", "00000000000110100110111101010011", "00000000001010011111011011101000", "00000000001101111100010000101011", "00000000010001011011101011011100", "00000000010100011101001100001110", "00000000010110110111111011010111", "00000000011001011100100011001110", "00000000011011000001000101000001", "00000000011011110110011001101011", "00000000011100110101011010101101", "00000000011100111000100111001001", "00000000011100000010010011110110", "00000000011011001100000001001001", "00000000011001101001110000001000", "00000000010111011110101111111000", "00000000010101011000011010110110", "00000000010010100101000110000100", "00000000001111001110100110101000", "00000000001011101000010001110010", "00000000000111101010110001101001", "00000000000011110111110111100001", "00000000000000000000001111000101", "11111111111100001000010110110010", "11111111111000010101011111010010", "11111111110100010111111111110011", "11111111110000110001101000001101", "11111111101101011011000110101000", "11111111101010100111101110111010", "11111111101000100001011000011101", "11111111100110010110011100011001", "11111111100100110100000000110101", "11111111100011111101101110100000", "11111111100011000111011001001111", "11111111100011001010100001111110", "11111111100100001001100001110000", "11111111100100111110110110111001", "11111111100110100011001110001010", "11111111101001000111111011100001", "11111111101011100010101010010000", "11111111101110100100000011000011", "11111111110010000011011110010011", "11111111110101100000010011100110", "11111111111001011000110011101110", "11111111111101001111110000101101", "00000000000001000110001100010011", "00000000000100111011010110101101", "00000000001000110110000100011000", "00000000001100100011001100111011", "00000000001111111100111100101110", "00000000010011011000011101001110", "00000000010110000010011101011010", "00000000011000001110011001100110", "00000000011010001001110001101111", "00000000011011101001100110111111", "00000000011100101111101100111100", "00000000011100111110111110110101", "00000000011100100010000101001000", "00000000011011101101011011000001", "00000000011010100101111101000001", "00000000011000110010100111000101", "00000000010110011000111000010000", "00000000010011101101110110100011", "00000000010000101000110111011000", "00000000001101001101010111100100", "00000000001001011000011111011000", "00000000000101100000000111110000", "00000000000001101011000011010010", "11111111111101110011001000100011", "11111111111001111101111100111010", "11111111110110000110001010001100", "11111111110010001111001000100111", "11111111101111001000001101110010", "11111111101100010010100101011110", "11111111101001001110010000101010", "11111111100111010011100111100001", "11111111100101011101100000111111", "11111111100011111011000101100000", "11111111100011100010000101111111", "11111111100011000001001110010100", "11111111100011100000010001001001", "11111111100100101110100010011001", "11111111100110001010011111010011", "11111111100111111101110110001011", "11111111101010001110100001001000", "11111111101101001111111110010101", "11111111110000001010100011011101", "11111111110011110110110101001001", "11111111110111100000101101001010", "11111111111011000110110011000111", "11111111111111100011100011101111", "00000000000011010000011011100001", "00000000000111000110111000010001", "00000000001011000101010001100010", "00000000001110100000100100111001", "00000000010001110111011001000101", "00000000010100011110101011001100", "00000000010111001010110100010001", "00000000011001100111100100010100", "00000000011010111000100111111110", "00000000011100001010011101001100", "00000000011101000000110101011111", "00000000011100110010110010100010", "00000000011100010001001110010001", "00000000011011001011101111101111", "00000000011001011000111110001100", "00000000010111010000110100101000", "00000000010100110000111100000000", "00000000010001111010110001010000", "00000000001110101001011001011111", "00000000001011001011110101100100", "00000000000111101111011111110100", "00000000000011110011100011001000", "11111111111111100000001111001010", "11111111111011100101111011111000", "11111111110111110000101110000110", "11111111110100000100010000100011", "11111111110000110001011000011001", "11111111101101010010110001011010", "11111111101010011010100000010111", "11111111101000010010001010010000", "11111111100110000101111110101010", "11111111100100011100011100011011", "11111111100011101100000001101011", "11111111100011011101011011110110", "11111111100011100010001100111110", "11111111100100000001100000101011", "11111111100101010001111110100001", "11111111100110111010001000111000", "11111111101001001010000110011111", "11111111101011111001001110100000", "11111111101110100000010111110100", "11111111110010001110100100101001", "11111111110101100011100011011010", "11111111111001010100001011010011", "11111111111101011100111011101011", "00000000000001000101001000100010", "00000000000101111011100111110111", "00000000001000111100010000101000", "00000000001101011001110110011011", "00000000010000100000110110000101", "00000000010011001110100011000111", "00000000010110111011000101001001", "00000000010111011000011100000011", "00000000011011111000001000001100", "00000000011010010100101101110110", "00000000011101111100000100110000", "00000000011101000001001111010011"));

end Outputs_test;

package body Outputs_Test is
end Outputs_Test;
