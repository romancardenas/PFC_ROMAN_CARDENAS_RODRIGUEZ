library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.ReSamplerTypes.all;

package CoeffConstants is

-- Declare constants

  constant coeffs : CoeffMatrix := 
  (
("000000000000000000",  "000000000000000000",  "000000000000000000",  "000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "000000000000000000",  "000000000000000000",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "000000000000000000",  "000000000000000000",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000000",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111011",  "000000000000111011",  "000000000000111011",  "000000000000111011",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111110",  "000000000000111110",  "000000000000111110",  "000000000000111110",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111110",  "000000000000111110",  "000000000000111110",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111011",  "000000000000111011",  "000000000000111011",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010100",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001110",  "000000000000001110",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001010",  "000000000000001010",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000110",  "000000000000000110",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000010",  "000000000000000010",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001100",  "111111111111001100",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001000",  "111111111111001000",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000100",  "111111111111000100",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111110",  "111111111110111110",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110110",  "111111111110110110",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110100",  "111111111110110100",  "111111111110110100",  "111111111110110011",  "111111111110110011",  "111111111110110011",  "111111111110110010",  "111111111110110010",  "111111111110110010",  "111111111110110001",  "111111111110110001",  "111111111110110001",  "111111111110110000",  "111111111110110000",  "111111111110110000",  "111111111110101111",  "111111111110101111",  "111111111110101111",  "111111111110101110",  "111111111110101110",  "111111111110101110",  "111111111110101101",  "111111111110101101",  "111111111110101101",  "111111111110101100",  "111111111110101100",  "111111111110101100",  "111111111110101011",  "111111111110101011",  "111111111110101011",  "111111111110101011",  "111111111110101010",  "111111111110101010",  "111111111110101010",  "111111111110101001",  "111111111110101001",  "111111111110101001",  "111111111110101000",  "111111111110101000",  "111111111110101000",  "111111111110100111",  "111111111110100111",  "111111111110100111",  "111111111110100110",  "111111111110100110",  "111111111110100110",  "111111111110100101",  "111111111110100101",  "111111111110100101",  "111111111110100100",  "111111111110100100",  "111111111110100100",  "111111111110100100",  "111111111110100011",  "111111111110100011",  "111111111110100011",  "111111111110100010",  "111111111110100010",  "111111111110100010",  "111111111110100001",  "111111111110100001",  "111111111110100001",  "111111111110100001",  "111111111110100000",  "111111111110100000",  "111111111110100000",  "111111111110011111",  "111111111110011111",  "111111111110011111",  "111111111110011110",  "111111111110011110",  "111111111110011110",  "111111111110011110",  "111111111110011101",  "111111111110011101",  "111111111110011101",  "111111111110011100",  "111111111110011100",  "111111111110011100",  "111111111110011011",  "111111111110011011",  "111111111110011011",  "111111111110011011",  "111111111110011010",  "111111111110011010",  "111111111110011010",  "111111111110011001",  "111111111110011001",  "111111111110011001",  "111111111110011001",  "111111111110011000",  "111111111110011000",  "111111111110011000",  "111111111110011000",  "111111111110010111",  "111111111110010111",  "111111111110010111",  "111111111110010110",  "111111111110010110",  "111111111110010110",  "111111111110010110",  "111111111110010101",  "111111111110010101",  "111111111110010101",  "111111111110010101",  "111111111110010100",  "111111111110010100",  "111111111110010100",  "111111111110010011",  "111111111110010011",  "111111111110010011",  "111111111110010011",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010001",  "111111111110010001",  "111111111110010001",  "111111111110010001",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110001110",  "111111111110001110",  "111111111110001110",  "111111111110001110",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001110",  "111111111110001110",  "111111111110001110",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110010001",  "111111111110010001",  "111111111110010001",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010011",  "111111111110010011",  "111111111110010011",  "111111111110010100",  "111111111110010100",  "111111111110010100",  "111111111110010100",  "111111111110010101",  "111111111110010101",  "111111111110010101",  "111111111110010110",  "111111111110010110",  "111111111110010110",  "111111111110010111",  "111111111110010111",  "111111111110010111",  "111111111110010111",  "111111111110011000",  "111111111110011000",  "111111111110011000",  "111111111110011001",  "111111111110011001",  "111111111110011001",  "111111111110011010",  "111111111110011010",  "111111111110011010",  "111111111110011011",  "111111111110011011",  "111111111110011011",  "111111111110011100",  "111111111110011100",  "111111111110011100",  "111111111110011101",  "111111111110011101",  "111111111110011101",  "111111111110011110",  "111111111110011110",  "111111111110011110",  "111111111110011111",  "111111111110011111",  "111111111110011111",  "111111111110100000",  "111111111110100000",  "111111111110100000",  "111111111110100001",  "111111111110100001",  "111111111110100001",  "111111111110100010",  "111111111110100010",  "111111111110100010",  "111111111110100011",  "111111111110100011",  "111111111110100011",  "111111111110100100",  "111111111110100100",  "111111111110100100",  "111111111110100101",  "111111111110100101",  "111111111110100101",  "111111111110100110",  "111111111110100110",  "111111111110100110",  "111111111110100111",  "111111111110100111",  "111111111110101000",  "111111111110101000",  "111111111110101000",  "111111111110101001",  "111111111110101001",  "111111111110101001",  "111111111110101010",  "111111111110101010",  "111111111110101010",  "111111111110101011",  "111111111110101011",  "111111111110101100",  "111111111110101100",  "111111111110101100",  "111111111110101101",  "111111111110101101",  "111111111110101101",  "111111111110101110",  "111111111110101110",  "111111111110101111",  "111111111110101111",  "111111111110101111",  "111111111110110000",  "111111111110110000",  "111111111110110001",  "111111111110110001",  "111111111110110001",  "111111111110110010",  "111111111110110010",  "111111111110110010",  "111111111110110011",  "111111111110110011",  "111111111110110100",  "111111111110110100",  "111111111110110100",  "111111111110110101",  "111111111110110101",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110111",  "111111111110110111",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111001",  "111111111110111001",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111011",  "111111111110111011",  "111111111110111100",  "111111111110111100",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111110",  "111111111110111110",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111111000000",  "111111111111000000",  "111111111111000001",  "111111111111000001",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000011",  "111111111111000011",  "111111111111000100",  "111111111111000100",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000110",  "111111111111000110",  "111111111111000111",  "111111111111000111",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001001",  "111111111111001001",  "111111111111001010",  "111111111111001010",  "111111111111001011",  "111111111111001011",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001101",  "111111111111001101",  "111111111111001110",  "111111111111001110",  "111111111111001111",  "111111111111001111",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111110",  "111111111111111111",  "111111111111111111"),("000000000000000000",  "000000000000000001",  "000000000000000001",  "000000000000000010",  "000000000000000010",  "000000000000000011",  "000000000000000011",  "000000000000000100",  "000000000000000100",  "000000000000000101",  "000000000000000101",  "000000000000000110",  "000000000000000110",  "000000000000000111",  "000000000000000111",  "000000000000001000",  "000000000000001000",  "000000000000001001",  "000000000000001001",  "000000000000001010",  "000000000000001010",  "000000000000001011",  "000000000000001011",  "000000000000001100",  "000000000000001100",  "000000000000001101",  "000000000000001101",  "000000000000001110",  "000000000000001110",  "000000000000001111",  "000000000000001111",  "000000000000010000",  "000000000000010000",  "000000000000010001",  "000000000000010001",  "000000000000010010",  "000000000000010010",  "000000000000010011",  "000000000000010011",  "000000000000010100",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010110",  "000000000000010111",  "000000000000010111",  "000000000000011000",  "000000000000011000",  "000000000000011001",  "000000000000011001",  "000000000000011010",  "000000000000011010",  "000000000000011011",  "000000000000011011",  "000000000000011100",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011110",  "000000000000011111",  "000000000000100000",  "000000000000100000",  "000000000000100001",  "000000000000100001",  "000000000000100010",  "000000000000100010",  "000000000000100011",  "000000000000100011",  "000000000000100100",  "000000000000100100",  "000000000000100101",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000100111",  "000000000000101000",  "000000000000101000",  "000000000000101001",  "000000000000101001",  "000000000000101010",  "000000000000101010",  "000000000000101011",  "000000000000101011",  "000000000000101100",  "000000000000101100",  "000000000000101101",  "000000000000101101",  "000000000000101110",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110000",  "000000000000110001",  "000000000000110001",  "000000000000110010",  "000000000000110010",  "000000000000110011",  "000000000000110011",  "000000000000110100",  "000000000000110100",  "000000000000110101",  "000000000000110101",  "000000000000110110",  "000000000000110110",  "000000000000110111",  "000000000000110111",  "000000000000111000",  "000000000000111000",  "000000000000111001",  "000000000000111010",  "000000000000111010",  "000000000000111011",  "000000000000111011",  "000000000000111100",  "000000000000111100",  "000000000000111101",  "000000000000111101",  "000000000000111110",  "000000000000111110",  "000000000000111111",  "000000000000111111",  "000000000001000000",  "000000000001000000",  "000000000001000001",  "000000000001000001",  "000000000001000010",  "000000000001000010",  "000000000001000011",  "000000000001000011",  "000000000001000100",  "000000000001000100",  "000000000001000101",  "000000000001000101",  "000000000001000110",  "000000000001000110",  "000000000001000111",  "000000000001000111",  "000000000001001000",  "000000000001001000",  "000000000001001001",  "000000000001001001",  "000000000001001010",  "000000000001001010",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001100",  "000000000001001100",  "000000000001001101",  "000000000001001101",  "000000000001001110",  "000000000001001110",  "000000000001001111",  "000000000001001111",  "000000000001010000",  "000000000001010000",  "000000000001010001",  "000000000001010001",  "000000000001010010",  "000000000001010010",  "000000000001010011",  "000000000001010011",  "000000000001010100",  "000000000001010100",  "000000000001010101",  "000000000001010101",  "000000000001010110",  "000000000001010110",  "000000000001010111",  "000000000001010111",  "000000000001011000",  "000000000001011000",  "000000000001011001",  "000000000001011001",  "000000000001011010",  "000000000001011010",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011100",  "000000000001011100",  "000000000001011101",  "000000000001011101",  "000000000001011110",  "000000000001011110",  "000000000001011111",  "000000000001011111",  "000000000001100000",  "000000000001100000",  "000000000001100001",  "000000000001100001",  "000000000001100010",  "000000000001100010",  "000000000001100011",  "000000000001100011",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100101",  "000000000001100101",  "000000000001100110",  "000000000001100110",  "000000000001100111",  "000000000001100111",  "000000000001101000",  "000000000001101000",  "000000000001101001",  "000000000001101001",  "000000000001101001",  "000000000001101010",  "000000000001101010",  "000000000001101011",  "000000000001101011",  "000000000001101100",  "000000000001101100",  "000000000001101101",  "000000000001101101",  "000000000001101110",  "000000000001101110",  "000000000001101110",  "000000000001101111",  "000000000001101111",  "000000000001110000",  "000000000001110000",  "000000000001110001",  "000000000001110001",  "000000000001110010",  "000000000001110010",  "000000000001110010",  "000000000001110011",  "000000000001110011",  "000000000001110100",  "000000000001110100",  "000000000001110101",  "000000000001110101",  "000000000001110110",  "000000000001110110",  "000000000001110110",  "000000000001110111",  "000000000001110111",  "000000000001111000",  "000000000001111000",  "000000000001111001",  "000000000001111001",  "000000000001111001",  "000000000001111010",  "000000000001111010",  "000000000001111011",  "000000000001111011",  "000000000001111100",  "000000000001111100",  "000000000001111100",  "000000000001111101",  "000000000001111101",  "000000000001111110",  "000000000001111110",  "000000000001111110",  "000000000001111111",  "000000000001111111",  "000000000010000000",  "000000000010000000",  "000000000010000001",  "000000000010000001",  "000000000010000001",  "000000000010000010",  "000000000010000010",  "000000000010000011",  "000000000010000011",  "000000000010000011",  "000000000010000100",  "000000000010000100",  "000000000010000101",  "000000000010000101",  "000000000010000101",  "000000000010000110",  "000000000010000110",  "000000000010000111",  "000000000010000111",  "000000000010000111",  "000000000010001000",  "000000000010001000",  "000000000010001001",  "000000000010001001",  "000000000010001001",  "000000000010001010",  "000000000010001010",  "000000000010001010",  "000000000010001011",  "000000000010001011",  "000000000010001100",  "000000000010001100",  "000000000010001100",  "000000000010001101",  "000000000010001101",  "000000000010001110",  "000000000010001110",  "000000000010001110",  "000000000010001111",  "000000000010001111",  "000000000010001111",  "000000000010010000",  "000000000010010000",  "000000000010010000",  "000000000010010001",  "000000000010010001",  "000000000010010010",  "000000000010010010",  "000000000010010010",  "000000000010010011",  "000000000010010011",  "000000000010010011",  "000000000010010100",  "000000000010010100",  "000000000010010100",  "000000000010010101",  "000000000010010101",  "000000000010010101",  "000000000010010110",  "000000000010010110",  "000000000010010111",  "000000000010010111",  "000000000010010111",  "000000000010011000",  "000000000010011000",  "000000000010011000",  "000000000010011001",  "000000000010011001",  "000000000010011001",  "000000000010011010",  "000000000010011010",  "000000000010011010",  "000000000010011011",  "000000000010011011",  "000000000010011011",  "000000000010011100",  "000000000010011100",  "000000000010011100",  "000000000010011101",  "000000000010011101",  "000000000010011101",  "000000000010011110",  "000000000010011110",  "000000000010011110",  "000000000010011110",  "000000000010011111",  "000000000010011111",  "000000000010011111",  "000000000010100000",  "000000000010100000",  "000000000010100000",  "000000000010100001",  "000000000010100001",  "000000000010100001",  "000000000010100010",  "000000000010100010",  "000000000010100010",  "000000000010100010",  "000000000010100011",  "000000000010100011",  "000000000010100011",  "000000000010100100",  "000000000010100100",  "000000000010100100",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100110",  "000000000010100110",  "000000000010100110",  "000000000010100111",  "000000000010100111",  "000000000010100111",  "000000000010100111",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010101001",  "000000000010101001",  "000000000010101001",  "000000000010101001",  "000000000010101010",  "000000000010101010",  "000000000010101010",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101010",  "000000000010101010",  "000000000010101010",  "000000000010101010",  "000000000010101001",  "000000000010101001",  "000000000010101001",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010100111",  "000000000010100111",  "000000000010100111",  "000000000010100110",  "000000000010100110",  "000000000010100110",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100100",  "000000000010100100",  "000000000010100100",  "000000000010100011",  "000000000010100011",  "000000000010100011",  "000000000010100010",  "000000000010100010",  "000000000010100010",  "000000000010100001",  "000000000010100001",  "000000000010100001",  "000000000010100000",  "000000000010100000",  "000000000010100000",  "000000000010011111",  "000000000010011111",  "000000000010011111",  "000000000010011110",  "000000000010011110",  "000000000010011110",  "000000000010011101",  "000000000010011101",  "000000000010011101",  "000000000010011100",  "000000000010011100",  "000000000010011100",  "000000000010011011",  "000000000010011011",  "000000000010011010",  "000000000010011010",  "000000000010011010",  "000000000010011001",  "000000000010011001",  "000000000010011001",  "000000000010011000",  "000000000010011000",  "000000000010011000",  "000000000010010111",  "000000000010010111",  "000000000010010110",  "000000000010010110",  "000000000010010110",  "000000000010010101",  "000000000010010101",  "000000000010010101",  "000000000010010100",  "000000000010010100",  "000000000010010011",  "000000000010010011",  "000000000010010011",  "000000000010010010",  "000000000010010010",  "000000000010010001",  "000000000010010001",  "000000000010010001",  "000000000010010000",  "000000000010010000",  "000000000010001111",  "000000000010001111",  "000000000010001111",  "000000000010001110",  "000000000010001110",  "000000000010001101",  "000000000010001101",  "000000000010001100",  "000000000010001100",  "000000000010001100",  "000000000010001011",  "000000000010001011",  "000000000010001010",  "000000000010001010",  "000000000010001001",  "000000000010001001",  "000000000010001001",  "000000000010001000",  "000000000010001000",  "000000000010000111",  "000000000010000111",  "000000000010000110",  "000000000010000110",  "000000000010000110",  "000000000010000101",  "000000000010000101",  "000000000010000100",  "000000000010000100",  "000000000010000011",  "000000000010000011",  "000000000010000010",  "000000000010000010",  "000000000010000010",  "000000000010000001",  "000000000010000001",  "000000000010000000",  "000000000010000000",  "000000000001111111",  "000000000001111111",  "000000000001111110",  "000000000001111110",  "000000000001111101",  "000000000001111101",  "000000000001111100",  "000000000001111100",  "000000000001111011",  "000000000001111011",  "000000000001111010",  "000000000001111010",  "000000000001111010",  "000000000001111001",  "000000000001111001",  "000000000001111000",  "000000000001111000",  "000000000001110111",  "000000000001110111",  "000000000001110110",  "000000000001110110",  "000000000001110101",  "000000000001110101",  "000000000001110100",  "000000000001110100",  "000000000001110011",  "000000000001110011",  "000000000001110010",  "000000000001110010",  "000000000001110001",  "000000000001110001",  "000000000001110000",  "000000000001110000",  "000000000001101111",  "000000000001101111",  "000000000001101110",  "000000000001101110",  "000000000001101101",  "000000000001101101",  "000000000001101100",  "000000000001101011",  "000000000001101011",  "000000000001101010",  "000000000001101010",  "000000000001101001",  "000000000001101001",  "000000000001101000",  "000000000001101000",  "000000000001100111",  "000000000001100111",  "000000000001100110",  "000000000001100110",  "000000000001100101",  "000000000001100101",  "000000000001100100",  "000000000001100100",  "000000000001100011",  "000000000001100010",  "000000000001100010",  "000000000001100001",  "000000000001100001",  "000000000001100000",  "000000000001100000",  "000000000001011111",  "000000000001011111",  "000000000001011110",  "000000000001011110",  "000000000001011101",  "000000000001011100",  "000000000001011100",  "000000000001011011",  "000000000001011011",  "000000000001011010",  "000000000001011010",  "000000000001011001",  "000000000001011001",  "000000000001011000",  "000000000001010111",  "000000000001010111",  "000000000001010110",  "000000000001010110",  "000000000001010101",  "000000000001010101",  "000000000001010100",  "000000000001010011",  "000000000001010011",  "000000000001010010",  "000000000001010010",  "000000000001010001",  "000000000001010001",  "000000000001010000",  "000000000001001111",  "000000000001001111",  "000000000001001110",  "000000000001001110",  "000000000001001101",  "000000000001001100",  "000000000001001100",  "000000000001001011",  "000000000001001011",  "000000000001001010",  "000000000001001010",  "000000000001001001",  "000000000001001000",  "000000000001001000",  "000000000001000111",  "000000000001000111",  "000000000001000110",  "000000000001000101",  "000000000001000101",  "000000000001000100",  "000000000001000100",  "000000000001000011",  "000000000001000010",  "000000000001000010",  "000000000001000001",  "000000000001000001",  "000000000001000000",  "000000000000111111",  "000000000000111111",  "000000000000111110",  "000000000000111101",  "000000000000111101",  "000000000000111100",  "000000000000111100",  "000000000000111011",  "000000000000111010",  "000000000000111010",  "000000000000111001",  "000000000000111001",  "000000000000111000",  "000000000000110111",  "000000000000110111",  "000000000000110110",  "000000000000110101",  "000000000000110101",  "000000000000110100",  "000000000000110100",  "000000000000110011",  "000000000000110010",  "000000000000110010",  "000000000000110001",  "000000000000110000",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101101",  "000000000000101101",  "000000000000101100",  "000000000000101011",  "000000000000101011",  "000000000000101010",  "000000000000101001",  "000000000000101001",  "000000000000101000",  "000000000000101000",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100100",  "000000000000100100",  "000000000000100011",  "000000000000100010",  "000000000000100010",  "000000000000100001",  "000000000000100000",  "000000000000100000",  "000000000000011111",  "000000000000011111",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011011",  "000000000000011011",  "000000000000011010",  "000000000000011001",  "000000000000011001",  "000000000000011000",  "000000000000010111",  "000000000000010111",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010011",  "000000000000010011",  "000000000000010010",  "000000000000010001",  "000000000000010001",  "000000000000010000",  "000000000000001111",  "000000000000001111",  "000000000000001110",  "000000000000001101",  "000000000000001101",  "000000000000001100",  "000000000000001011",  "000000000000001011",  "000000000000001010",  "000000000000001001",  "000000000000001001",  "000000000000001000",  "000000000000000111",  "000000000000000111",  "000000000000000110",  "000000000000000101",  "000000000000000101",  "000000000000000100",  "000000000000000011",  "000000000000000011",  "000000000000000010",  "000000000000000001",  "000000000000000001"),("000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111001111",  "111111111111001110",  "111111111111001110",  "111111111111001101",  "111111111111001100",  "111111111111001011",  "111111111111001011",  "111111111111001010",  "111111111111001001",  "111111111111001001",  "111111111111001000",  "111111111111000111",  "111111111111000111",  "111111111111000110",  "111111111111000101",  "111111111111000101",  "111111111111000100",  "111111111111000011",  "111111111111000011",  "111111111111000010",  "111111111111000001",  "111111111111000001",  "111111111111000000",  "111111111110111111",  "111111111110111111",  "111111111110111110",  "111111111110111101",  "111111111110111100",  "111111111110111100",  "111111111110111011",  "111111111110111010",  "111111111110111010",  "111111111110111001",  "111111111110111000",  "111111111110111000",  "111111111110110111",  "111111111110110110",  "111111111110110110",  "111111111110110101",  "111111111110110100",  "111111111110110100",  "111111111110110011",  "111111111110110010",  "111111111110110010",  "111111111110110001",  "111111111110110000",  "111111111110110000",  "111111111110101111",  "111111111110101110",  "111111111110101110",  "111111111110101101",  "111111111110101100",  "111111111110101100",  "111111111110101011",  "111111111110101010",  "111111111110101010",  "111111111110101001",  "111111111110101000",  "111111111110101000",  "111111111110100111",  "111111111110100110",  "111111111110100110",  "111111111110100101",  "111111111110100100",  "111111111110100100",  "111111111110100011",  "111111111110100010",  "111111111110100010",  "111111111110100001",  "111111111110100000",  "111111111110100000",  "111111111110011111",  "111111111110011110",  "111111111110011110",  "111111111110011101",  "111111111110011100",  "111111111110011100",  "111111111110011011",  "111111111110011010",  "111111111110011010",  "111111111110011001",  "111111111110011000",  "111111111110011000",  "111111111110010111",  "111111111110010110",  "111111111110010110",  "111111111110010101",  "111111111110010100",  "111111111110010100",  "111111111110010011",  "111111111110010010",  "111111111110010010",  "111111111110010001",  "111111111110010001",  "111111111110010000",  "111111111110001111",  "111111111110001111",  "111111111110001110",  "111111111110001101",  "111111111110001101",  "111111111110001100",  "111111111110001011",  "111111111110001011",  "111111111110001010",  "111111111110001001",  "111111111110001001",  "111111111110001000",  "111111111110001000",  "111111111110000111",  "111111111110000110",  "111111111110000110",  "111111111110000101",  "111111111110000100",  "111111111110000100",  "111111111110000011",  "111111111110000010",  "111111111110000010",  "111111111110000001",  "111111111110000001",  "111111111110000000",  "111111111101111111",  "111111111101111111",  "111111111101111110",  "111111111101111101",  "111111111101111101",  "111111111101111100",  "111111111101111100",  "111111111101111011",  "111111111101111010",  "111111111101111010",  "111111111101111001",  "111111111101111000",  "111111111101111000",  "111111111101110111",  "111111111101110111",  "111111111101110110",  "111111111101110101",  "111111111101110101",  "111111111101110100",  "111111111101110100",  "111111111101110011",  "111111111101110010",  "111111111101110010",  "111111111101110001",  "111111111101110001",  "111111111101110000",  "111111111101101111",  "111111111101101111",  "111111111101101110",  "111111111101101110",  "111111111101101101",  "111111111101101100",  "111111111101101100",  "111111111101101011",  "111111111101101011",  "111111111101101010",  "111111111101101001",  "111111111101101001",  "111111111101101000",  "111111111101101000",  "111111111101100111",  "111111111101100110",  "111111111101100110",  "111111111101100101",  "111111111101100101",  "111111111101100100",  "111111111101100100",  "111111111101100011",  "111111111101100010",  "111111111101100010",  "111111111101100001",  "111111111101100001",  "111111111101100000",  "111111111101100000",  "111111111101011111",  "111111111101011110",  "111111111101011110",  "111111111101011101",  "111111111101011101",  "111111111101011100",  "111111111101011100",  "111111111101011011",  "111111111101011010",  "111111111101011010",  "111111111101011001",  "111111111101011001",  "111111111101011000",  "111111111101011000",  "111111111101010111",  "111111111101010111",  "111111111101010110",  "111111111101010101",  "111111111101010101",  "111111111101010100",  "111111111101010100",  "111111111101010011",  "111111111101010011",  "111111111101010010",  "111111111101010010",  "111111111101010001",  "111111111101010001",  "111111111101010000",  "111111111101001111",  "111111111101001111",  "111111111101001110",  "111111111101001110",  "111111111101001101",  "111111111101001101",  "111111111101001100",  "111111111101001100",  "111111111101001011",  "111111111101001011",  "111111111101001010",  "111111111101001010",  "111111111101001001",  "111111111101001001",  "111111111101001000",  "111111111101001000",  "111111111101000111",  "111111111101000111",  "111111111101000110",  "111111111101000110",  "111111111101000101",  "111111111101000101",  "111111111101000100",  "111111111101000100",  "111111111101000011",  "111111111101000011",  "111111111101000010",  "111111111101000010",  "111111111101000001",  "111111111101000001",  "111111111101000000",  "111111111101000000",  "111111111100111111",  "111111111100111111",  "111111111100111110",  "111111111100111110",  "111111111100111101",  "111111111100111101",  "111111111100111100",  "111111111100111100",  "111111111100111011",  "111111111100111011",  "111111111100111010",  "111111111100111010",  "111111111100111001",  "111111111100111001",  "111111111100111001",  "111111111100111000",  "111111111100111000",  "111111111100110111",  "111111111100110111",  "111111111100110110",  "111111111100110110",  "111111111100110101",  "111111111100110101",  "111111111100110100",  "111111111100110100",  "111111111100110100",  "111111111100110011",  "111111111100110011",  "111111111100110010",  "111111111100110010",  "111111111100110001",  "111111111100110001",  "111111111100110000",  "111111111100110000",  "111111111100110000",  "111111111100101111",  "111111111100101111",  "111111111100101110",  "111111111100101110",  "111111111100101101",  "111111111100101101",  "111111111100101101",  "111111111100101100",  "111111111100101100",  "111111111100101011",  "111111111100101011",  "111111111100101011",  "111111111100101010",  "111111111100101010",  "111111111100101001",  "111111111100101001",  "111111111100101001",  "111111111100101000",  "111111111100101000",  "111111111100100111",  "111111111100100111",  "111111111100100111",  "111111111100100110",  "111111111100100110",  "111111111100100101",  "111111111100100101",  "111111111100100101",  "111111111100100100",  "111111111100100100",  "111111111100100100",  "111111111100100011",  "111111111100100011",  "111111111100100010",  "111111111100100010",  "111111111100100010",  "111111111100100001",  "111111111100100001",  "111111111100100001",  "111111111100100000",  "111111111100100000",  "111111111100100000",  "111111111100011111",  "111111111100011111",  "111111111100011110",  "111111111100011110",  "111111111100011110",  "111111111100011101",  "111111111100011101",  "111111111100011101",  "111111111100011100",  "111111111100011100",  "111111111100011100",  "111111111100011011",  "111111111100011011",  "111111111100011011",  "111111111100011010",  "111111111100011010",  "111111111100011010",  "111111111100011001",  "111111111100011001",  "111111111100011001",  "111111111100011001",  "111111111100011000",  "111111111100011000",  "111111111100011000",  "111111111100010111",  "111111111100010111",  "111111111100010111",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010101",  "111111111100010101",  "111111111100010101",  "111111111100010100",  "111111111100010100",  "111111111100010100",  "111111111100010100",  "111111111100010011",  "111111111100010011",  "111111111100010011",  "111111111100010010",  "111111111100010010",  "111111111100010010",  "111111111100010010",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010010",  "111111111100010010",  "111111111100010010",  "111111111100010011",  "111111111100010011",  "111111111100010011",  "111111111100010011",  "111111111100010100",  "111111111100010100",  "111111111100010100",  "111111111100010101",  "111111111100010101",  "111111111100010101",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010111",  "111111111100010111",  "111111111100010111",  "111111111100011000",  "111111111100011000",  "111111111100011000",  "111111111100011001",  "111111111100011001",  "111111111100011001",  "111111111100011010",  "111111111100011010",  "111111111100011010",  "111111111100011011",  "111111111100011011",  "111111111100011011",  "111111111100011100",  "111111111100011100",  "111111111100011100",  "111111111100011101",  "111111111100011101",  "111111111100011110",  "111111111100011110",  "111111111100011110",  "111111111100011111",  "111111111100011111",  "111111111100011111",  "111111111100100000",  "111111111100100000",  "111111111100100000",  "111111111100100001",  "111111111100100001",  "111111111100100010",  "111111111100100010",  "111111111100100010",  "111111111100100011",  "111111111100100011",  "111111111100100100",  "111111111100100100",  "111111111100100100",  "111111111100100101",  "111111111100100101",  "111111111100100110",  "111111111100100110",  "111111111100100110",  "111111111100100111",  "111111111100100111",  "111111111100101000",  "111111111100101000",  "111111111100101001",  "111111111100101001",  "111111111100101001",  "111111111100101010",  "111111111100101010",  "111111111100101011",  "111111111100101011",  "111111111100101100",  "111111111100101100",  "111111111100101101",  "111111111100101101",  "111111111100101101",  "111111111100101110",  "111111111100101110",  "111111111100101111",  "111111111100101111",  "111111111100110000",  "111111111100110000",  "111111111100110001",  "111111111100110001",  "111111111100110010",  "111111111100110010",  "111111111100110011",  "111111111100110011",  "111111111100110011",  "111111111100110100",  "111111111100110100",  "111111111100110101",  "111111111100110101",  "111111111100110110",  "111111111100110110",  "111111111100110111",  "111111111100110111",  "111111111100111000",  "111111111100111000",  "111111111100111001",  "111111111100111001",  "111111111100111010",  "111111111100111010",  "111111111100111011",  "111111111100111011",  "111111111100111100",  "111111111100111100",  "111111111100111101",  "111111111100111110",  "111111111100111110",  "111111111100111111",  "111111111100111111",  "111111111101000000",  "111111111101000000",  "111111111101000001",  "111111111101000001",  "111111111101000010",  "111111111101000010",  "111111111101000011",  "111111111101000011",  "111111111101000100",  "111111111101000100",  "111111111101000101",  "111111111101000110",  "111111111101000110",  "111111111101000111",  "111111111101000111",  "111111111101001000",  "111111111101001000",  "111111111101001001",  "111111111101001010",  "111111111101001010",  "111111111101001011",  "111111111101001011",  "111111111101001100",  "111111111101001100",  "111111111101001101",  "111111111101001110",  "111111111101001110",  "111111111101001111",  "111111111101001111",  "111111111101010000",  "111111111101010001",  "111111111101010001",  "111111111101010010",  "111111111101010010",  "111111111101010011",  "111111111101010100",  "111111111101010100",  "111111111101010101",  "111111111101010101",  "111111111101010110",  "111111111101010111",  "111111111101010111",  "111111111101011000",  "111111111101011000",  "111111111101011001",  "111111111101011010",  "111111111101011010",  "111111111101011011",  "111111111101011100",  "111111111101011100",  "111111111101011101",  "111111111101011101",  "111111111101011110",  "111111111101011111",  "111111111101011111",  "111111111101100000",  "111111111101100001",  "111111111101100001",  "111111111101100010",  "111111111101100011",  "111111111101100011",  "111111111101100100",  "111111111101100100",  "111111111101100101",  "111111111101100110",  "111111111101100110",  "111111111101100111",  "111111111101101000",  "111111111101101000",  "111111111101101001",  "111111111101101010",  "111111111101101010",  "111111111101101011",  "111111111101101100",  "111111111101101100",  "111111111101101101",  "111111111101101110",  "111111111101101111",  "111111111101101111",  "111111111101110000",  "111111111101110001",  "111111111101110001",  "111111111101110010",  "111111111101110011",  "111111111101110011",  "111111111101110100",  "111111111101110101",  "111111111101110101",  "111111111101110110",  "111111111101110111",  "111111111101111000",  "111111111101111000",  "111111111101111001",  "111111111101111010",  "111111111101111010",  "111111111101111011",  "111111111101111100",  "111111111101111100",  "111111111101111101",  "111111111101111110",  "111111111101111111",  "111111111101111111",  "111111111110000000",  "111111111110000001",  "111111111110000010",  "111111111110000010",  "111111111110000011",  "111111111110000100",  "111111111110000100",  "111111111110000101",  "111111111110000110",  "111111111110000111",  "111111111110000111",  "111111111110001000",  "111111111110001001",  "111111111110001010",  "111111111110001010",  "111111111110001011",  "111111111110001100",  "111111111110001101",  "111111111110001101",  "111111111110001110",  "111111111110001111",  "111111111110010000",  "111111111110010000",  "111111111110010001",  "111111111110010010",  "111111111110010011",  "111111111110010011",  "111111111110010100",  "111111111110010101",  "111111111110010110",  "111111111110010110",  "111111111110010111",  "111111111110011000",  "111111111110011001",  "111111111110011010",  "111111111110011010",  "111111111110011011",  "111111111110011100",  "111111111110011101",  "111111111110011101",  "111111111110011110",  "111111111110011111",  "111111111110100000",  "111111111110100001",  "111111111110100001",  "111111111110100010",  "111111111110100011",  "111111111110100100",  "111111111110100100",  "111111111110100101",  "111111111110100110",  "111111111110100111",  "111111111110101000",  "111111111110101000",  "111111111110101001",  "111111111110101010",  "111111111110101011",  "111111111110101100",  "111111111110101100",  "111111111110101101",  "111111111110101110",  "111111111110101111",  "111111111110110000",  "111111111110110001",  "111111111110110001",  "111111111110110010",  "111111111110110011",  "111111111110110100",  "111111111110110101",  "111111111110110101",  "111111111110110110",  "111111111110110111",  "111111111110111000",  "111111111110111001",  "111111111110111001",  "111111111110111010",  "111111111110111011",  "111111111110111100",  "111111111110111101",  "111111111110111110",  "111111111110111110",  "111111111110111111",  "111111111111000000",  "111111111111000001",  "111111111111000010",  "111111111111000011",  "111111111111000011",  "111111111111000100",  "111111111111000101",  "111111111111000110",  "111111111111000111",  "111111111111001000",  "111111111111001000",  "111111111111001001",  "111111111111001010",  "111111111111001011",  "111111111111001100",  "111111111111001101",  "111111111111001110",  "111111111111001110",  "111111111111001111",  "111111111111010000",  "111111111111010001",  "111111111111010010",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010110",  "111111111111010111",  "111111111111011000",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011100",  "111111111111011101",  "111111111111011110",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100010",  "111111111111100011",  "111111111111100100",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111101000",  "111111111111101001",  "111111111111101010",  "111111111111101011",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101111",  "111111111111110000",  "111111111111110001",  "111111111111110010",  "111111111111110011",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110111",  "111111111111111000",  "111111111111111001",  "111111111111111010",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111110",  "111111111111111111"),("000000000000000000",  "000000000000000001",  "000000000000000010",  "000000000000000011",  "000000000000000100",  "000000000000000100",  "000000000000000101",  "000000000000000110",  "000000000000000111",  "000000000000001000",  "000000000000001001",  "000000000000001010",  "000000000000001011",  "000000000000001100",  "000000000000001100",  "000000000000001101",  "000000000000001110",  "000000000000001111",  "000000000000010000",  "000000000000010001",  "000000000000010010",  "000000000000010011",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010111",  "000000000000011000",  "000000000000011001",  "000000000000011010",  "000000000000011011",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011111",  "000000000000100000",  "000000000000100001",  "000000000000100010",  "000000000000100011",  "000000000000100100",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000101000",  "000000000000101001",  "000000000000101010",  "000000000000101011",  "000000000000101100",  "000000000000101101",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110001",  "000000000000110010",  "000000000000110011",  "000000000000110100",  "000000000000110101",  "000000000000110110",  "000000000000110111",  "000000000000111000",  "000000000000111000",  "000000000000111001",  "000000000000111010",  "000000000000111011",  "000000000000111100",  "000000000000111101",  "000000000000111110",  "000000000000111111",  "000000000001000000",  "000000000001000001",  "000000000001000001",  "000000000001000010",  "000000000001000011",  "000000000001000100",  "000000000001000101",  "000000000001000110",  "000000000001000111",  "000000000001001000",  "000000000001001001",  "000000000001001010",  "000000000001001010",  "000000000001001011",  "000000000001001100",  "000000000001001101",  "000000000001001110",  "000000000001001111",  "000000000001010000",  "000000000001010001",  "000000000001010010",  "000000000001010011",  "000000000001010011",  "000000000001010100",  "000000000001010101",  "000000000001010110",  "000000000001010111",  "000000000001011000",  "000000000001011001",  "000000000001011010",  "000000000001011011",  "000000000001011011",  "000000000001011100",  "000000000001011101",  "000000000001011110",  "000000000001011111",  "000000000001100000",  "000000000001100001",  "000000000001100010",  "000000000001100011",  "000000000001100011",  "000000000001100100",  "000000000001100101",  "000000000001100110",  "000000000001100111",  "000000000001101000",  "000000000001101001",  "000000000001101010",  "000000000001101011",  "000000000001101011",  "000000000001101100",  "000000000001101101",  "000000000001101110",  "000000000001101111",  "000000000001110000",  "000000000001110001",  "000000000001110010",  "000000000001110010",  "000000000001110011",  "000000000001110100",  "000000000001110101",  "000000000001110110",  "000000000001110111",  "000000000001111000",  "000000000001111001",  "000000000001111001",  "000000000001111010",  "000000000001111011",  "000000000001111100",  "000000000001111101",  "000000000001111110",  "000000000001111111",  "000000000010000000",  "000000000010000000",  "000000000010000001",  "000000000010000010",  "000000000010000011",  "000000000010000100",  "000000000010000101",  "000000000010000110",  "000000000010000110",  "000000000010000111",  "000000000010001000",  "000000000010001001",  "000000000010001010",  "000000000010001011",  "000000000010001100",  "000000000010001100",  "000000000010001101",  "000000000010001110",  "000000000010001111",  "000000000010010000",  "000000000010010001",  "000000000010010010",  "000000000010010010",  "000000000010010011",  "000000000010010100",  "000000000010010101",  "000000000010010110",  "000000000010010111",  "000000000010010111",  "000000000010011000",  "000000000010011001",  "000000000010011010",  "000000000010011011",  "000000000010011100",  "000000000010011101",  "000000000010011101",  "000000000010011110",  "000000000010011111",  "000000000010100000",  "000000000010100001",  "000000000010100010",  "000000000010100010",  "000000000010100011",  "000000000010100100",  "000000000010100101",  "000000000010100110",  "000000000010100110",  "000000000010100111",  "000000000010101000",  "000000000010101001",  "000000000010101010",  "000000000010101011",  "000000000010101011",  "000000000010101100",  "000000000010101101",  "000000000010101110",  "000000000010101111",  "000000000010101111",  "000000000010110000",  "000000000010110001",  "000000000010110010",  "000000000010110011",  "000000000010110011",  "000000000010110100",  "000000000010110101",  "000000000010110110",  "000000000010110111",  "000000000010110111",  "000000000010111000",  "000000000010111001",  "000000000010111010",  "000000000010111011",  "000000000010111011",  "000000000010111100",  "000000000010111101",  "000000000010111110",  "000000000010111111",  "000000000010111111",  "000000000011000000",  "000000000011000001",  "000000000011000010",  "000000000011000011",  "000000000011000011",  "000000000011000100",  "000000000011000101",  "000000000011000110",  "000000000011000110",  "000000000011000111",  "000000000011001000",  "000000000011001001",  "000000000011001001",  "000000000011001010",  "000000000011001011",  "000000000011001100",  "000000000011001100",  "000000000011001101",  "000000000011001110",  "000000000011001111",  "000000000011010000",  "000000000011010000",  "000000000011010001",  "000000000011010010",  "000000000011010010",  "000000000011010011",  "000000000011010100",  "000000000011010101",  "000000000011010101",  "000000000011010110",  "000000000011010111",  "000000000011011000",  "000000000011011000",  "000000000011011001",  "000000000011011010",  "000000000011011011",  "000000000011011011",  "000000000011011100",  "000000000011011101",  "000000000011011101",  "000000000011011110",  "000000000011011111",  "000000000011100000",  "000000000011100000",  "000000000011100001",  "000000000011100010",  "000000000011100010",  "000000000011100011",  "000000000011100100",  "000000000011100101",  "000000000011100101",  "000000000011100110",  "000000000011100111",  "000000000011100111",  "000000000011101000",  "000000000011101001",  "000000000011101001",  "000000000011101010",  "000000000011101011",  "000000000011101100",  "000000000011101100",  "000000000011101101",  "000000000011101110",  "000000000011101110",  "000000000011101111",  "000000000011110000",  "000000000011110000",  "000000000011110001",  "000000000011110010",  "000000000011110010",  "000000000011110011",  "000000000011110100",  "000000000011110100",  "000000000011110101",  "000000000011110110",  "000000000011110110",  "000000000011110111",  "000000000011111000",  "000000000011111000",  "000000000011111001",  "000000000011111001",  "000000000011111010",  "000000000011111011",  "000000000011111011",  "000000000011111100",  "000000000011111101",  "000000000011111101",  "000000000011111110",  "000000000011111111",  "000000000011111111",  "000000000100000000",  "000000000100000000",  "000000000100000001",  "000000000100000010",  "000000000100000010",  "000000000100000011",  "000000000100000011",  "000000000100000100",  "000000000100000101",  "000000000100000101",  "000000000100000110",  "000000000100000110",  "000000000100000111",  "000000000100001000",  "000000000100001000",  "000000000100001001",  "000000000100001001",  "000000000100001010",  "000000000100001011",  "000000000100001011",  "000000000100001100",  "000000000100001100",  "000000000100001101",  "000000000100001101",  "000000000100001110",  "000000000100001111",  "000000000100001111",  "000000000100010000",  "000000000100010000",  "000000000100010001",  "000000000100010001",  "000000000100010010",  "000000000100010011",  "000000000100010011",  "000000000100010100",  "000000000100010100",  "000000000100010101",  "000000000100010101",  "000000000100010110",  "000000000100010110",  "000000000100010111",  "000000000100010111",  "000000000100011000",  "000000000100011000",  "000000000100011001",  "000000000100011001",  "000000000100011010",  "000000000100011011",  "000000000100011011",  "000000000100011100",  "000000000100011100",  "000000000100011101",  "000000000100011101",  "000000000100011110",  "000000000100011110",  "000000000100011111",  "000000000100011111",  "000000000100100000",  "000000000100100000",  "000000000100100001",  "000000000100100001",  "000000000100100001",  "000000000100100010",  "000000000100100010",  "000000000100100011",  "000000000100100011",  "000000000100100100",  "000000000100100100",  "000000000100100101",  "000000000100100101",  "000000000100100110",  "000000000100100110",  "000000000100100111",  "000000000100100111",  "000000000100101000",  "000000000100101000",  "000000000100101000",  "000000000100101001",  "000000000100101001",  "000000000100101010",  "000000000100101010",  "000000000100101011",  "000000000100101011",  "000000000100101011",  "000000000100101100",  "000000000100101100",  "000000000100101101",  "000000000100101101",  "000000000100101110",  "000000000100101110",  "000000000100101110",  "000000000100101111",  "000000000100101111",  "000000000100110000",  "000000000100110000",  "000000000100110000",  "000000000100110001",  "000000000100110001",  "000000000100110010",  "000000000100110010",  "000000000100110010",  "000000000100110011",  "000000000100110011",  "000000000100110011",  "000000000100110100",  "000000000100110100",  "000000000100110100",  "000000000100110101",  "000000000100110101",  "000000000100110110",  "000000000100110110",  "000000000100110110",  "000000000100110111",  "000000000100110111",  "000000000100110111",  "000000000100111000",  "000000000100111000",  "000000000100111000",  "000000000100111001",  "000000000100111001",  "000000000100111001",  "000000000100111010",  "000000000100111010",  "000000000100111010",  "000000000100111011",  "000000000100111011",  "000000000100111011",  "000000000100111011",  "000000000100111100",  "000000000100111100",  "000000000100111100",  "000000000100111101",  "000000000100111101",  "000000000100111101",  "000000000100111110",  "000000000100111110",  "000000000100111110",  "000000000100111110",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000101000000",  "000000000101000000",  "000000000101000000",  "000000000101000000",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000000",  "000000000101000000",  "000000000101000000",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000100111110",  "000000000100111110",  "000000000100111110",  "000000000100111101",  "000000000100111101",  "000000000100111101",  "000000000100111101",  "000000000100111100",  "000000000100111100",  "000000000100111100",  "000000000100111011",  "000000000100111011",  "000000000100111011",  "000000000100111010",  "000000000100111010",  "000000000100111010",  "000000000100111001",  "000000000100111001",  "000000000100111001",  "000000000100111000",  "000000000100111000",  "000000000100111000",  "000000000100110111",  "000000000100110111",  "000000000100110111",  "000000000100110110",  "000000000100110110",  "000000000100110110",  "000000000100110101",  "000000000100110101",  "000000000100110100",  "000000000100110100",  "000000000100110100",  "000000000100110011",  "000000000100110011",  "000000000100110011",  "000000000100110010",  "000000000100110010",  "000000000100110001",  "000000000100110001",  "000000000100110001",  "000000000100110000",  "000000000100110000",  "000000000100101111",  "000000000100101111",  "000000000100101110",  "000000000100101110",  "000000000100101110",  "000000000100101101",  "000000000100101101",  "000000000100101100",  "000000000100101100",  "000000000100101011",  "000000000100101011",  "000000000100101010",  "000000000100101010",  "000000000100101010",  "000000000100101001",  "000000000100101001",  "000000000100101000",  "000000000100101000",  "000000000100100111",  "000000000100100111",  "000000000100100110",  "000000000100100110",  "000000000100100101",  "000000000100100101",  "000000000100100100",  "000000000100100100",  "000000000100100011",  "000000000100100011",  "000000000100100010",  "000000000100100010",  "000000000100100001",  "000000000100100001",  "000000000100100000",  "000000000100100000",  "000000000100011111",  "000000000100011111",  "000000000100011110",  "000000000100011110",  "000000000100011101",  "000000000100011101",  "000000000100011100",  "000000000100011100",  "000000000100011011",  "000000000100011010",  "000000000100011010",  "000000000100011001",  "000000000100011001",  "000000000100011000",  "000000000100011000",  "000000000100010111",  "000000000100010111",  "000000000100010110",  "000000000100010101",  "000000000100010101",  "000000000100010100",  "000000000100010100",  "000000000100010011",  "000000000100010011",  "000000000100010010",  "000000000100010001",  "000000000100010001",  "000000000100010000",  "000000000100010000",  "000000000100001111",  "000000000100001110",  "000000000100001110",  "000000000100001101",  "000000000100001100",  "000000000100001100",  "000000000100001011",  "000000000100001011",  "000000000100001010",  "000000000100001001",  "000000000100001001",  "000000000100001000",  "000000000100000111",  "000000000100000111",  "000000000100000110",  "000000000100000110",  "000000000100000101",  "000000000100000100",  "000000000100000100",  "000000000100000011",  "000000000100000010",  "000000000100000010",  "000000000100000001",  "000000000100000000",  "000000000100000000",  "000000000011111111",  "000000000011111110",  "000000000011111110",  "000000000011111101",  "000000000011111100",  "000000000011111011",  "000000000011111011",  "000000000011111010",  "000000000011111001",  "000000000011111001",  "000000000011111000",  "000000000011110111",  "000000000011110111",  "000000000011110110",  "000000000011110101",  "000000000011110100",  "000000000011110100",  "000000000011110011",  "000000000011110010",  "000000000011110010",  "000000000011110001",  "000000000011110000",  "000000000011101111",  "000000000011101111",  "000000000011101110",  "000000000011101101",  "000000000011101100",  "000000000011101100",  "000000000011101011",  "000000000011101010",  "000000000011101001",  "000000000011101001",  "000000000011101000",  "000000000011100111",  "000000000011100110",  "000000000011100110",  "000000000011100101",  "000000000011100100",  "000000000011100011",  "000000000011100010",  "000000000011100010",  "000000000011100001",  "000000000011100000",  "000000000011011111",  "000000000011011111",  "000000000011011110",  "000000000011011101",  "000000000011011100",  "000000000011011011",  "000000000011011011",  "000000000011011010",  "000000000011011001",  "000000000011011000",  "000000000011010111",  "000000000011010110",  "000000000011010110",  "000000000011010101",  "000000000011010100",  "000000000011010011",  "000000000011010010",  "000000000011010010",  "000000000011010001",  "000000000011010000",  "000000000011001111",  "000000000011001110",  "000000000011001101",  "000000000011001100",  "000000000011001100",  "000000000011001011",  "000000000011001010",  "000000000011001001",  "000000000011001000",  "000000000011000111",  "000000000011000111",  "000000000011000110",  "000000000011000101",  "000000000011000100",  "000000000011000011",  "000000000011000010",  "000000000011000001",  "000000000011000000",  "000000000011000000",  "000000000010111111",  "000000000010111110",  "000000000010111101",  "000000000010111100",  "000000000010111011",  "000000000010111010",  "000000000010111001",  "000000000010111000",  "000000000010111000",  "000000000010110111",  "000000000010110110",  "000000000010110101",  "000000000010110100",  "000000000010110011",  "000000000010110010",  "000000000010110001",  "000000000010110000",  "000000000010101111",  "000000000010101110",  "000000000010101101",  "000000000010101101",  "000000000010101100",  "000000000010101011",  "000000000010101010",  "000000000010101001",  "000000000010101000",  "000000000010100111",  "000000000010100110",  "000000000010100101",  "000000000010100100",  "000000000010100011",  "000000000010100010",  "000000000010100001",  "000000000010100000",  "000000000010011111",  "000000000010011110",  "000000000010011101",  "000000000010011101",  "000000000010011100",  "000000000010011011",  "000000000010011010",  "000000000010011001",  "000000000010011000",  "000000000010010111",  "000000000010010110",  "000000000010010101",  "000000000010010100",  "000000000010010011",  "000000000010010010",  "000000000010010001",  "000000000010010000",  "000000000010001111",  "000000000010001110",  "000000000010001101",  "000000000010001100",  "000000000010001011",  "000000000010001010",  "000000000010001001",  "000000000010001000",  "000000000010000111",  "000000000010000110",  "000000000010000101",  "000000000010000100",  "000000000010000011",  "000000000010000010",  "000000000010000001",  "000000000010000000",  "000000000001111111",  "000000000001111110",  "000000000001111101",  "000000000001111100",  "000000000001111011",  "000000000001111010",  "000000000001111001",  "000000000001111000",  "000000000001110111",  "000000000001110110",  "000000000001110101",  "000000000001110100",  "000000000001110011",  "000000000001110001",  "000000000001110000",  "000000000001101111",  "000000000001101110",  "000000000001101101",  "000000000001101100",  "000000000001101011",  "000000000001101010",  "000000000001101001",  "000000000001101000",  "000000000001100111",  "000000000001100110",  "000000000001100101",  "000000000001100100",  "000000000001100011",  "000000000001100010",  "000000000001100001",  "000000000001100000",  "000000000001011111",  "000000000001011110",  "000000000001011100",  "000000000001011011",  "000000000001011010",  "000000000001011001",  "000000000001011000",  "000000000001010111",  "000000000001010110",  "000000000001010101",  "000000000001010100",  "000000000001010011",  "000000000001010010",  "000000000001010001",  "000000000001010000",  "000000000001001110",  "000000000001001101",  "000000000001001100",  "000000000001001011",  "000000000001001010",  "000000000001001001",  "000000000001001000",  "000000000001000111",  "000000000001000110",  "000000000001000101",  "000000000001000100",  "000000000001000010",  "000000000001000001",  "000000000001000000",  "000000000000111111",  "000000000000111110",  "000000000000111101",  "000000000000111100",  "000000000000111011",  "000000000000111010",  "000000000000111001",  "000000000000110111",  "000000000000110110",  "000000000000110101",  "000000000000110100",  "000000000000110011",  "000000000000110010",  "000000000000110001",  "000000000000110000",  "000000000000101111",  "000000000000101101",  "000000000000101100",  "000000000000101011",  "000000000000101010",  "000000000000101001",  "000000000000101000",  "000000000000100111",  "000000000000100110",  "000000000000100100",  "000000000000100011",  "000000000000100010",  "000000000000100001",  "000000000000100000",  "000000000000011111",  "000000000000011110",  "000000000000011101",  "000000000000011011",  "000000000000011010",  "000000000000011001",  "000000000000011000",  "000000000000010111",  "000000000000010110",  "000000000000010101",  "000000000000010011",  "000000000000010010",  "000000000000010001",  "000000000000010000",  "000000000000001111",  "000000000000001110",  "000000000000001101",  "000000000000001011",  "000000000000001010",  "000000000000001001",  "000000000000001000",  "000000000000000111",  "000000000000000110",  "000000000000000101",  "000000000000000011",  "000000000000000010",  "000000000000000001"),("000000000000000000",  "111111111111111111",  "111111111111111110",  "111111111111111101",  "111111111111111011",  "111111111111111010",  "111111111111111001",  "111111111111111000",  "111111111111110111",  "111111111111110110",  "111111111111110100",  "111111111111110011",  "111111111111110010",  "111111111111110001",  "111111111111110000",  "111111111111101111",  "111111111111101110",  "111111111111101100",  "111111111111101011",  "111111111111101010",  "111111111111101001",  "111111111111101000",  "111111111111100111",  "111111111111100101",  "111111111111100100",  "111111111111100011",  "111111111111100010",  "111111111111100001",  "111111111111100000",  "111111111111011110",  "111111111111011101",  "111111111111011100",  "111111111111011011",  "111111111111011010",  "111111111111011001",  "111111111111011000",  "111111111111010110",  "111111111111010101",  "111111111111010100",  "111111111111010011",  "111111111111010010",  "111111111111010001",  "111111111111001111",  "111111111111001110",  "111111111111001101",  "111111111111001100",  "111111111111001011",  "111111111111001010",  "111111111111001000",  "111111111111000111",  "111111111111000110",  "111111111111000101",  "111111111111000100",  "111111111111000011",  "111111111111000001",  "111111111111000000",  "111111111110111111",  "111111111110111110",  "111111111110111101",  "111111111110111100",  "111111111110111010",  "111111111110111001",  "111111111110111000",  "111111111110110111",  "111111111110110110",  "111111111110110101",  "111111111110110011",  "111111111110110010",  "111111111110110001",  "111111111110110000",  "111111111110101111",  "111111111110101110",  "111111111110101100",  "111111111110101011",  "111111111110101010",  "111111111110101001",  "111111111110101000",  "111111111110100111",  "111111111110100110",  "111111111110100100",  "111111111110100011",  "111111111110100010",  "111111111110100001",  "111111111110100000",  "111111111110011111",  "111111111110011101",  "111111111110011100",  "111111111110011011",  "111111111110011010",  "111111111110011001",  "111111111110011000",  "111111111110010110",  "111111111110010101",  "111111111110010100",  "111111111110010011",  "111111111110010010",  "111111111110010001",  "111111111110010000",  "111111111110001110",  "111111111110001101",  "111111111110001100",  "111111111110001011",  "111111111110001010",  "111111111110001001",  "111111111110001000",  "111111111110000110",  "111111111110000101",  "111111111110000100",  "111111111110000011",  "111111111110000010",  "111111111110000001",  "111111111101111111",  "111111111101111110",  "111111111101111101",  "111111111101111100",  "111111111101111011",  "111111111101111010",  "111111111101111001",  "111111111101110111",  "111111111101110110",  "111111111101110101",  "111111111101110100",  "111111111101110011",  "111111111101110010",  "111111111101110001",  "111111111101110000",  "111111111101101110",  "111111111101101101",  "111111111101101100",  "111111111101101011",  "111111111101101010",  "111111111101101001",  "111111111101101000",  "111111111101100110",  "111111111101100101",  "111111111101100100",  "111111111101100011",  "111111111101100010",  "111111111101100001",  "111111111101100000",  "111111111101011111",  "111111111101011110",  "111111111101011100",  "111111111101011011",  "111111111101011010",  "111111111101011001",  "111111111101011000",  "111111111101010111",  "111111111101010110",  "111111111101010101",  "111111111101010011",  "111111111101010010",  "111111111101010001",  "111111111101010000",  "111111111101001111",  "111111111101001110",  "111111111101001101",  "111111111101001100",  "111111111101001011",  "111111111101001010",  "111111111101001000",  "111111111101000111",  "111111111101000110",  "111111111101000101",  "111111111101000100",  "111111111101000011",  "111111111101000010",  "111111111101000001",  "111111111101000000",  "111111111100111111",  "111111111100111110",  "111111111100111100",  "111111111100111011",  "111111111100111010",  "111111111100111001",  "111111111100111000",  "111111111100110111",  "111111111100110110",  "111111111100110101",  "111111111100110100",  "111111111100110011",  "111111111100110010",  "111111111100110001",  "111111111100110000",  "111111111100101110",  "111111111100101101",  "111111111100101100",  "111111111100101011",  "111111111100101010",  "111111111100101001",  "111111111100101000",  "111111111100100111",  "111111111100100110",  "111111111100100101",  "111111111100100100",  "111111111100100011",  "111111111100100010",  "111111111100100001",  "111111111100100000",  "111111111100011111",  "111111111100011110",  "111111111100011101",  "111111111100011100",  "111111111100011011",  "111111111100011001",  "111111111100011000",  "111111111100010111",  "111111111100010110",  "111111111100010101",  "111111111100010100",  "111111111100010011",  "111111111100010010",  "111111111100010001",  "111111111100010000",  "111111111100001111",  "111111111100001110",  "111111111100001101",  "111111111100001100",  "111111111100001011",  "111111111100001010",  "111111111100001001",  "111111111100001000",  "111111111100000111",  "111111111100000110",  "111111111100000101",  "111111111100000100",  "111111111100000011",  "111111111100000010",  "111111111100000001",  "111111111100000000",  "111111111011111111",  "111111111011111110",  "111111111011111101",  "111111111011111100",  "111111111011111011",  "111111111011111010",  "111111111011111001",  "111111111011111000",  "111111111011110111",  "111111111011110110",  "111111111011110101",  "111111111011110100",  "111111111011110011",  "111111111011110011",  "111111111011110010",  "111111111011110001",  "111111111011110000",  "111111111011101111",  "111111111011101110",  "111111111011101101",  "111111111011101100",  "111111111011101011",  "111111111011101010",  "111111111011101001",  "111111111011101000",  "111111111011100111",  "111111111011100110",  "111111111011100101",  "111111111011100100",  "111111111011100011",  "111111111011100011",  "111111111011100010",  "111111111011100001",  "111111111011100000",  "111111111011011111",  "111111111011011110",  "111111111011011101",  "111111111011011100",  "111111111011011011",  "111111111011011010",  "111111111011011001",  "111111111011011001",  "111111111011011000",  "111111111011010111",  "111111111011010110",  "111111111011010101",  "111111111011010100",  "111111111011010011",  "111111111011010010",  "111111111011010001",  "111111111011010001",  "111111111011010000",  "111111111011001111",  "111111111011001110",  "111111111011001101",  "111111111011001100",  "111111111011001011",  "111111111011001010",  "111111111011001010",  "111111111011001001",  "111111111011001000",  "111111111011000111",  "111111111011000110",  "111111111011000101",  "111111111011000101",  "111111111011000100",  "111111111011000011",  "111111111011000010",  "111111111011000001",  "111111111011000000",  "111111111011000000",  "111111111010111111",  "111111111010111110",  "111111111010111101",  "111111111010111100",  "111111111010111011",  "111111111010111011",  "111111111010111010",  "111111111010111001",  "111111111010111000",  "111111111010110111",  "111111111010110111",  "111111111010110110",  "111111111010110101",  "111111111010110100",  "111111111010110011",  "111111111010110011",  "111111111010110010",  "111111111010110001",  "111111111010110000",  "111111111010110000",  "111111111010101111",  "111111111010101110",  "111111111010101101",  "111111111010101100",  "111111111010101100",  "111111111010101011",  "111111111010101010",  "111111111010101001",  "111111111010101001",  "111111111010101000",  "111111111010100111",  "111111111010100111",  "111111111010100110",  "111111111010100101",  "111111111010100100",  "111111111010100100",  "111111111010100011",  "111111111010100010",  "111111111010100001",  "111111111010100001",  "111111111010100000",  "111111111010011111",  "111111111010011111",  "111111111010011110",  "111111111010011101",  "111111111010011101",  "111111111010011100",  "111111111010011011",  "111111111010011010",  "111111111010011010",  "111111111010011001",  "111111111010011000",  "111111111010011000",  "111111111010010111",  "111111111010010110",  "111111111010010110",  "111111111010010101",  "111111111010010100",  "111111111010010100",  "111111111010010011",  "111111111010010010",  "111111111010010010",  "111111111010010001",  "111111111010010001",  "111111111010010000",  "111111111010001111",  "111111111010001111",  "111111111010001110",  "111111111010001101",  "111111111010001101",  "111111111010001100",  "111111111010001100",  "111111111010001011",  "111111111010001010",  "111111111010001010",  "111111111010001001",  "111111111010001000",  "111111111010001000",  "111111111010000111",  "111111111010000111",  "111111111010000110",  "111111111010000110",  "111111111010000101",  "111111111010000100",  "111111111010000100",  "111111111010000011",  "111111111010000011",  "111111111010000010",  "111111111010000010",  "111111111010000001",  "111111111010000000",  "111111111010000000",  "111111111001111111",  "111111111001111111",  "111111111001111110",  "111111111001111110",  "111111111001111101",  "111111111001111101",  "111111111001111100",  "111111111001111100",  "111111111001111011",  "111111111001111011",  "111111111001111010",  "111111111001111010",  "111111111001111001",  "111111111001111001",  "111111111001111000",  "111111111001111000",  "111111111001110111",  "111111111001110111",  "111111111001110110",  "111111111001110110",  "111111111001110101",  "111111111001110101",  "111111111001110100",  "111111111001110100",  "111111111001110011",  "111111111001110011",  "111111111001110010",  "111111111001110010",  "111111111001110010",  "111111111001110001",  "111111111001110001",  "111111111001110000",  "111111111001110000",  "111111111001101111",  "111111111001101111",  "111111111001101111",  "111111111001101110",  "111111111001101110",  "111111111001101101",  "111111111001101101",  "111111111001101100",  "111111111001101100",  "111111111001101100",  "111111111001101011",  "111111111001101011",  "111111111001101010",  "111111111001101010",  "111111111001101010",  "111111111001101001",  "111111111001101001",  "111111111001101001",  "111111111001101000",  "111111111001101000",  "111111111001101000",  "111111111001100111",  "111111111001100111",  "111111111001100110",  "111111111001100110",  "111111111001100110",  "111111111001100101",  "111111111001100101",  "111111111001100101",  "111111111001100101",  "111111111001100100",  "111111111001100100",  "111111111001100100",  "111111111001100011",  "111111111001100011",  "111111111001100011",  "111111111001100010",  "111111111001100010",  "111111111001100010",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100000",  "111111111001100000",  "111111111001100000",  "111111111001100000",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001100000",  "111111111001100000",  "111111111001100000",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100010",  "111111111001100010",  "111111111001100010",  "111111111001100011",  "111111111001100011",  "111111111001100011",  "111111111001100100",  "111111111001100100",  "111111111001100100",  "111111111001100100",  "111111111001100101",  "111111111001100101",  "111111111001100110",  "111111111001100110",  "111111111001100110",  "111111111001100111",  "111111111001100111",  "111111111001100111",  "111111111001101000",  "111111111001101000",  "111111111001101000",  "111111111001101001",  "111111111001101001",  "111111111001101010",  "111111111001101010",  "111111111001101010",  "111111111001101011",  "111111111001101011",  "111111111001101011",  "111111111001101100",  "111111111001101100",  "111111111001101101",  "111111111001101101",  "111111111001101110",  "111111111001101110",  "111111111001101110",  "111111111001101111",  "111111111001101111",  "111111111001110000",  "111111111001110000",  "111111111001110001",  "111111111001110001",  "111111111001110010",  "111111111001110010",  "111111111001110010",  "111111111001110011",  "111111111001110011",  "111111111001110100",  "111111111001110100",  "111111111001110101",  "111111111001110101",  "111111111001110110",  "111111111001110110",  "111111111001110111",  "111111111001110111",  "111111111001111000",  "111111111001111000",  "111111111001111001",  "111111111001111001",  "111111111001111010",  "111111111001111011",  "111111111001111011",  "111111111001111100",  "111111111001111100",  "111111111001111101",  "111111111001111101",  "111111111001111110",  "111111111001111110",  "111111111001111111",  "111111111001111111",  "111111111010000000",  "111111111010000001",  "111111111010000001",  "111111111010000010",  "111111111010000010",  "111111111010000011",  "111111111010000100",  "111111111010000100",  "111111111010000101",  "111111111010000101",  "111111111010000110",  "111111111010000111",  "111111111010000111",  "111111111010001000",  "111111111010001000",  "111111111010001001",  "111111111010001010",  "111111111010001010",  "111111111010001011",  "111111111010001100",  "111111111010001100",  "111111111010001101",  "111111111010001110",  "111111111010001110",  "111111111010001111",  "111111111010010000",  "111111111010010000",  "111111111010010001",  "111111111010010010",  "111111111010010010",  "111111111010010011",  "111111111010010100",  "111111111010010100",  "111111111010010101",  "111111111010010110",  "111111111010010110",  "111111111010010111",  "111111111010011000",  "111111111010011001",  "111111111010011001",  "111111111010011010",  "111111111010011011",  "111111111010011011",  "111111111010011100",  "111111111010011101",  "111111111010011110",  "111111111010011110",  "111111111010011111",  "111111111010100000",  "111111111010100001",  "111111111010100001",  "111111111010100010",  "111111111010100011",  "111111111010100100",  "111111111010100101",  "111111111010100101",  "111111111010100110",  "111111111010100111",  "111111111010101000",  "111111111010101000",  "111111111010101001",  "111111111010101010",  "111111111010101011",  "111111111010101100",  "111111111010101101",  "111111111010101101",  "111111111010101110",  "111111111010101111",  "111111111010110000",  "111111111010110001",  "111111111010110001",  "111111111010110010",  "111111111010110011",  "111111111010110100",  "111111111010110101",  "111111111010110110",  "111111111010110111",  "111111111010110111",  "111111111010111000",  "111111111010111001",  "111111111010111010",  "111111111010111011",  "111111111010111100",  "111111111010111101",  "111111111010111101",  "111111111010111110",  "111111111010111111",  "111111111011000000",  "111111111011000001",  "111111111011000010",  "111111111011000011",  "111111111011000100",  "111111111011000101",  "111111111011000110",  "111111111011000111",  "111111111011000111",  "111111111011001000",  "111111111011001001",  "111111111011001010",  "111111111011001011",  "111111111011001100",  "111111111011001101",  "111111111011001110",  "111111111011001111",  "111111111011010000",  "111111111011010001",  "111111111011010010",  "111111111011010011",  "111111111011010100",  "111111111011010101",  "111111111011010110",  "111111111011010111",  "111111111011011000",  "111111111011011001",  "111111111011011010",  "111111111011011011",  "111111111011011100",  "111111111011011101",  "111111111011011110",  "111111111011011111",  "111111111011100000",  "111111111011100001",  "111111111011100010",  "111111111011100011",  "111111111011100100",  "111111111011100101",  "111111111011100110",  "111111111011100111",  "111111111011101000",  "111111111011101001",  "111111111011101010",  "111111111011101011",  "111111111011101100",  "111111111011101101",  "111111111011101110",  "111111111011101111",  "111111111011110000",  "111111111011110001",  "111111111011110010",  "111111111011110011",  "111111111011110100",  "111111111011110101",  "111111111011110110",  "111111111011110111",  "111111111011111001",  "111111111011111010",  "111111111011111011",  "111111111011111100",  "111111111011111101",  "111111111011111110",  "111111111011111111",  "111111111100000000",  "111111111100000001",  "111111111100000010",  "111111111100000011",  "111111111100000101",  "111111111100000110",  "111111111100000111",  "111111111100001000",  "111111111100001001",  "111111111100001010",  "111111111100001011",  "111111111100001100",  "111111111100001110",  "111111111100001111",  "111111111100010000",  "111111111100010001",  "111111111100010010",  "111111111100010011",  "111111111100010100",  "111111111100010110",  "111111111100010111",  "111111111100011000",  "111111111100011001",  "111111111100011010",  "111111111100011011",  "111111111100011101",  "111111111100011110",  "111111111100011111",  "111111111100100000",  "111111111100100001",  "111111111100100010",  "111111111100100100",  "111111111100100101",  "111111111100100110",  "111111111100100111",  "111111111100101000",  "111111111100101010",  "111111111100101011",  "111111111100101100",  "111111111100101101",  "111111111100101110",  "111111111100110000",  "111111111100110001",  "111111111100110010",  "111111111100110011",  "111111111100110100",  "111111111100110110",  "111111111100110111",  "111111111100111000",  "111111111100111001",  "111111111100111011",  "111111111100111100",  "111111111100111101",  "111111111100111110",  "111111111101000000",  "111111111101000001",  "111111111101000010",  "111111111101000011",  "111111111101000101",  "111111111101000110",  "111111111101000111",  "111111111101001000",  "111111111101001010",  "111111111101001011",  "111111111101001100",  "111111111101001101",  "111111111101001111",  "111111111101010000",  "111111111101010001",  "111111111101010011",  "111111111101010100",  "111111111101010101",  "111111111101010110",  "111111111101011000",  "111111111101011001",  "111111111101011010",  "111111111101011100",  "111111111101011101",  "111111111101011110",  "111111111101011111",  "111111111101100001",  "111111111101100010",  "111111111101100011",  "111111111101100101",  "111111111101100110",  "111111111101100111",  "111111111101101001",  "111111111101101010",  "111111111101101011",  "111111111101101101",  "111111111101101110",  "111111111101101111",  "111111111101110001",  "111111111101110010",  "111111111101110011",  "111111111101110100",  "111111111101110110",  "111111111101110111",  "111111111101111001",  "111111111101111010",  "111111111101111011",  "111111111101111101",  "111111111101111110",  "111111111101111111",  "111111111110000001",  "111111111110000010",  "111111111110000011",  "111111111110000101",  "111111111110000110",  "111111111110000111",  "111111111110001001",  "111111111110001010",  "111111111110001011",  "111111111110001101",  "111111111110001110",  "111111111110010000",  "111111111110010001",  "111111111110010010",  "111111111110010100",  "111111111110010101",  "111111111110010110",  "111111111110011000",  "111111111110011001",  "111111111110011011",  "111111111110011100",  "111111111110011101",  "111111111110011111",  "111111111110100000",  "111111111110100001",  "111111111110100011",  "111111111110100100",  "111111111110100110",  "111111111110100111",  "111111111110101000",  "111111111110101010",  "111111111110101011",  "111111111110101101",  "111111111110101110",  "111111111110101111",  "111111111110110001",  "111111111110110010",  "111111111110110100",  "111111111110110101",  "111111111110110111",  "111111111110111000",  "111111111110111001",  "111111111110111011",  "111111111110111100",  "111111111110111110",  "111111111110111111",  "111111111111000000",  "111111111111000010",  "111111111111000011",  "111111111111000101",  "111111111111000110",  "111111111111001000",  "111111111111001001",  "111111111111001010",  "111111111111001100",  "111111111111001101",  "111111111111001111",  "111111111111010000",  "111111111111010010",  "111111111111010011",  "111111111111010100",  "111111111111010110",  "111111111111010111",  "111111111111011001",  "111111111111011010",  "111111111111011100",  "111111111111011101",  "111111111111011111",  "111111111111100000",  "111111111111100001",  "111111111111100011",  "111111111111100100",  "111111111111100110",  "111111111111100111",  "111111111111101001",  "111111111111101010",  "111111111111101100",  "111111111111101101",  "111111111111101110",  "111111111111110000",  "111111111111110001",  "111111111111110011",  "111111111111110100",  "111111111111110110",  "111111111111110111",  "111111111111111001",  "111111111111111010",  "111111111111111100",  "111111111111111101",  "111111111111111111"),("000000000000000000",  "000000000000000001",  "000000000000000011",  "000000000000000100",  "000000000000000110",  "000000000000000111",  "000000000000001001",  "000000000000001010",  "000000000000001100",  "000000000000001101",  "000000000000001111",  "000000000000010000",  "000000000000010010",  "000000000000010011",  "000000000000010101",  "000000000000010110",  "000000000000011000",  "000000000000011001",  "000000000000011010",  "000000000000011100",  "000000000000011101",  "000000000000011111",  "000000000000100000",  "000000000000100010",  "000000000000100011",  "000000000000100101",  "000000000000100110",  "000000000000101000",  "000000000000101001",  "000000000000101011",  "000000000000101100",  "000000000000101110",  "000000000000101111",  "000000000000110001",  "000000000000110010",  "000000000000110100",  "000000000000110101",  "000000000000110111",  "000000000000111000",  "000000000000111001",  "000000000000111011",  "000000000000111100",  "000000000000111110",  "000000000000111111",  "000000000001000001",  "000000000001000010",  "000000000001000100",  "000000000001000101",  "000000000001000111",  "000000000001001000",  "000000000001001010",  "000000000001001011",  "000000000001001101",  "000000000001001110",  "000000000001010000",  "000000000001010001",  "000000000001010011",  "000000000001010100",  "000000000001010110",  "000000000001010111",  "000000000001011001",  "000000000001011010",  "000000000001011100",  "000000000001011101",  "000000000001011110",  "000000000001100000",  "000000000001100001",  "000000000001100011",  "000000000001100100",  "000000000001100110",  "000000000001100111",  "000000000001101001",  "000000000001101010",  "000000000001101100",  "000000000001101101",  "000000000001101111",  "000000000001110000",  "000000000001110010",  "000000000001110011",  "000000000001110101",  "000000000001110110",  "000000000001111000",  "000000000001111001",  "000000000001111011",  "000000000001111100",  "000000000001111101",  "000000000001111111",  "000000000010000000",  "000000000010000010",  "000000000010000011",  "000000000010000101",  "000000000010000110",  "000000000010001000",  "000000000010001001",  "000000000010001011",  "000000000010001100",  "000000000010001110",  "000000000010001111",  "000000000010010001",  "000000000010010010",  "000000000010010011",  "000000000010010101",  "000000000010010110",  "000000000010011000",  "000000000010011001",  "000000000010011011",  "000000000010011100",  "000000000010011110",  "000000000010011111",  "000000000010100001",  "000000000010100010",  "000000000010100011",  "000000000010100101",  "000000000010100110",  "000000000010101000",  "000000000010101001",  "000000000010101011",  "000000000010101100",  "000000000010101110",  "000000000010101111",  "000000000010110001",  "000000000010110010",  "000000000010110011",  "000000000010110101",  "000000000010110110",  "000000000010111000",  "000000000010111001",  "000000000010111011",  "000000000010111100",  "000000000010111101",  "000000000010111111",  "000000000011000000",  "000000000011000010",  "000000000011000011",  "000000000011000101",  "000000000011000110",  "000000000011000111",  "000000000011001001",  "000000000011001010",  "000000000011001100",  "000000000011001101",  "000000000011001111",  "000000000011010000",  "000000000011010001",  "000000000011010011",  "000000000011010100",  "000000000011010110",  "000000000011010111",  "000000000011011001",  "000000000011011010",  "000000000011011011",  "000000000011011101",  "000000000011011110",  "000000000011100000",  "000000000011100001",  "000000000011100010",  "000000000011100100",  "000000000011100101",  "000000000011100111",  "000000000011101000",  "000000000011101001",  "000000000011101011",  "000000000011101100",  "000000000011101110",  "000000000011101111",  "000000000011110000",  "000000000011110010",  "000000000011110011",  "000000000011110100",  "000000000011110110",  "000000000011110111",  "000000000011111001",  "000000000011111010",  "000000000011111011",  "000000000011111101",  "000000000011111110",  "000000000011111111",  "000000000100000001",  "000000000100000010",  "000000000100000011",  "000000000100000101",  "000000000100000110",  "000000000100001000",  "000000000100001001",  "000000000100001010",  "000000000100001100",  "000000000100001101",  "000000000100001110",  "000000000100010000",  "000000000100010001",  "000000000100010010",  "000000000100010100",  "000000000100010101",  "000000000100010110",  "000000000100011000",  "000000000100011001",  "000000000100011010",  "000000000100011100",  "000000000100011101",  "000000000100011110",  "000000000100100000",  "000000000100100001",  "000000000100100010",  "000000000100100100",  "000000000100100101",  "000000000100100110",  "000000000100100111",  "000000000100101001",  "000000000100101010",  "000000000100101011",  "000000000100101101",  "000000000100101110",  "000000000100101111",  "000000000100110001",  "000000000100110010",  "000000000100110011",  "000000000100110100",  "000000000100110110",  "000000000100110111",  "000000000100111000",  "000000000100111010",  "000000000100111011",  "000000000100111100",  "000000000100111101",  "000000000100111111",  "000000000101000000",  "000000000101000001",  "000000000101000010",  "000000000101000100",  "000000000101000101",  "000000000101000110",  "000000000101000111",  "000000000101001001",  "000000000101001010",  "000000000101001011",  "000000000101001100",  "000000000101001110",  "000000000101001111",  "000000000101010000",  "000000000101010001",  "000000000101010011",  "000000000101010100",  "000000000101010101",  "000000000101010110",  "000000000101010111",  "000000000101011001",  "000000000101011010",  "000000000101011011",  "000000000101011100",  "000000000101011101",  "000000000101011111",  "000000000101100000",  "000000000101100001",  "000000000101100010",  "000000000101100011",  "000000000101100101",  "000000000101100110",  "000000000101100111",  "000000000101101000",  "000000000101101001",  "000000000101101010",  "000000000101101100",  "000000000101101101",  "000000000101101110",  "000000000101101111",  "000000000101110000",  "000000000101110001",  "000000000101110011",  "000000000101110100",  "000000000101110101",  "000000000101110110",  "000000000101110111",  "000000000101111000",  "000000000101111001",  "000000000101111010",  "000000000101111100",  "000000000101111101",  "000000000101111110",  "000000000101111111",  "000000000110000000",  "000000000110000001",  "000000000110000010",  "000000000110000011",  "000000000110000100",  "000000000110000110",  "000000000110000111",  "000000000110001000",  "000000000110001001",  "000000000110001010",  "000000000110001011",  "000000000110001100",  "000000000110001101",  "000000000110001110",  "000000000110001111",  "000000000110010000",  "000000000110010001",  "000000000110010010",  "000000000110010011",  "000000000110010101",  "000000000110010110",  "000000000110010111",  "000000000110011000",  "000000000110011001",  "000000000110011010",  "000000000110011011",  "000000000110011100",  "000000000110011101",  "000000000110011110",  "000000000110011111",  "000000000110100000",  "000000000110100001",  "000000000110100010",  "000000000110100011",  "000000000110100100",  "000000000110100101",  "000000000110100110",  "000000000110100111",  "000000000110101000",  "000000000110101001",  "000000000110101010",  "000000000110101011",  "000000000110101100",  "000000000110101101",  "000000000110101110",  "000000000110101111",  "000000000110110000",  "000000000110110001",  "000000000110110001",  "000000000110110010",  "000000000110110011",  "000000000110110100",  "000000000110110101",  "000000000110110110",  "000000000110110111",  "000000000110111000",  "000000000110111001",  "000000000110111010",  "000000000110111011",  "000000000110111100",  "000000000110111101",  "000000000110111101",  "000000000110111110",  "000000000110111111",  "000000000111000000",  "000000000111000001",  "000000000111000010",  "000000000111000011",  "000000000111000100",  "000000000111000101",  "000000000111000101",  "000000000111000110",  "000000000111000111",  "000000000111001000",  "000000000111001001",  "000000000111001010",  "000000000111001010",  "000000000111001011",  "000000000111001100",  "000000000111001101",  "000000000111001110",  "000000000111001111",  "000000000111001111",  "000000000111010000",  "000000000111010001",  "000000000111010010",  "000000000111010011",  "000000000111010011",  "000000000111010100",  "000000000111010101",  "000000000111010110",  "000000000111010111",  "000000000111010111",  "000000000111011000",  "000000000111011001",  "000000000111011010",  "000000000111011010",  "000000000111011011",  "000000000111011100",  "000000000111011101",  "000000000111011101",  "000000000111011110",  "000000000111011111",  "000000000111100000",  "000000000111100000",  "000000000111100001",  "000000000111100010",  "000000000111100011",  "000000000111100011",  "000000000111100100",  "000000000111100101",  "000000000111100101",  "000000000111100110",  "000000000111100111",  "000000000111100111",  "000000000111101000",  "000000000111101001",  "000000000111101001",  "000000000111101010",  "000000000111101011",  "000000000111101011",  "000000000111101100",  "000000000111101101",  "000000000111101101",  "000000000111101110",  "000000000111101111",  "000000000111101111",  "000000000111110000",  "000000000111110000",  "000000000111110001",  "000000000111110010",  "000000000111110010",  "000000000111110011",  "000000000111110100",  "000000000111110100",  "000000000111110101",  "000000000111110101",  "000000000111110110",  "000000000111110110",  "000000000111110111",  "000000000111111000",  "000000000111111000",  "000000000111111001",  "000000000111111001",  "000000000111111010",  "000000000111111010",  "000000000111111011",  "000000000111111011",  "000000000111111100",  "000000000111111101",  "000000000111111101",  "000000000111111110",  "000000000111111110",  "000000000111111111",  "000000000111111111",  "000000001000000000",  "000000001000000000",  "000000001000000001",  "000000001000000001",  "000000001000000010",  "000000001000000010",  "000000001000000010",  "000000001000000011",  "000000001000000011",  "000000001000000100",  "000000001000000100",  "000000001000000101",  "000000001000000101",  "000000001000000110",  "000000001000000110",  "000000001000000111",  "000000001000000111",  "000000001000000111",  "000000001000001000",  "000000001000001000",  "000000001000001001",  "000000001000001001",  "000000001000001001",  "000000001000001010",  "000000001000001010",  "000000001000001011",  "000000001000001011",  "000000001000001011",  "000000001000001100",  "000000001000001100",  "000000001000001100",  "000000001000001101",  "000000001000001101",  "000000001000001101",  "000000001000001110",  "000000001000001110",  "000000001000001110",  "000000001000001111",  "000000001000001111",  "000000001000001111",  "000000001000010000",  "000000001000010000",  "000000001000010000",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010010",  "000000001000010010",  "000000001000010010",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010010",  "000000001000010010",  "000000001000010010",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010000",  "000000001000010000",  "000000001000010000",  "000000001000001111",  "000000001000001111",  "000000001000001111",  "000000001000001110",  "000000001000001110",  "000000001000001110",  "000000001000001101",  "000000001000001101",  "000000001000001101",  "000000001000001100",  "000000001000001100",  "000000001000001011",  "000000001000001011",  "000000001000001011",  "000000001000001010",  "000000001000001010",  "000000001000001010",  "000000001000001001",  "000000001000001001",  "000000001000001000",  "000000001000001000",  "000000001000000111",  "000000001000000111",  "000000001000000111",  "000000001000000110",  "000000001000000110",  "000000001000000101",  "000000001000000101",  "000000001000000100",  "000000001000000100",  "000000001000000011",  "000000001000000011",  "000000001000000010",  "000000001000000010",  "000000001000000001",  "000000001000000001",  "000000001000000000",  "000000001000000000",  "000000000111111111",  "000000000111111111",  "000000000111111110",  "000000000111111110",  "000000000111111101",  "000000000111111101",  "000000000111111100",  "000000000111111100",  "000000000111111011",  "000000000111111011",  "000000000111111010",  "000000000111111010",  "000000000111111001",  "000000000111111000",  "000000000111111000",  "000000000111110111",  "000000000111110111",  "000000000111110110",  "000000000111110101",  "000000000111110101",  "000000000111110100",  "000000000111110100",  "000000000111110011",  "000000000111110010",  "000000000111110010",  "000000000111110001",  "000000000111110000",  "000000000111110000",  "000000000111101111",  "000000000111101110",  "000000000111101110",  "000000000111101101",  "000000000111101100",  "000000000111101100",  "000000000111101011",  "000000000111101010",  "000000000111101010",  "000000000111101001",  "000000000111101000",  "000000000111101000",  "000000000111100111",  "000000000111100110",  "000000000111100101",  "000000000111100101",  "000000000111100100",  "000000000111100011",  "000000000111100011",  "000000000111100010",  "000000000111100001",  "000000000111100000",  "000000000111011111",  "000000000111011111",  "000000000111011110",  "000000000111011101",  "000000000111011100",  "000000000111011100",  "000000000111011011",  "000000000111011010",  "000000000111011001",  "000000000111011000",  "000000000111011000",  "000000000111010111",  "000000000111010110",  "000000000111010101",  "000000000111010100",  "000000000111010011",  "000000000111010011",  "000000000111010010",  "000000000111010001",  "000000000111010000",  "000000000111001111",  "000000000111001110",  "000000000111001110",  "000000000111001101",  "000000000111001100",  "000000000111001011",  "000000000111001010",  "000000000111001001",  "000000000111001000",  "000000000111000111",  "000000000111000110",  "000000000111000110",  "000000000111000101",  "000000000111000100",  "000000000111000011",  "000000000111000010",  "000000000111000001",  "000000000111000000",  "000000000110111111",  "000000000110111110",  "000000000110111101",  "000000000110111100",  "000000000110111011",  "000000000110111010",  "000000000110111001",  "000000000110111000",  "000000000110110111",  "000000000110110110",  "000000000110110101",  "000000000110110100",  "000000000110110011",  "000000000110110010",  "000000000110110001",  "000000000110110000",  "000000000110101111",  "000000000110101110",  "000000000110101101",  "000000000110101100",  "000000000110101011",  "000000000110101010",  "000000000110101001",  "000000000110101000",  "000000000110100111",  "000000000110100110",  "000000000110100101",  "000000000110100100",  "000000000110100011",  "000000000110100010",  "000000000110100001",  "000000000110100000",  "000000000110011110",  "000000000110011101",  "000000000110011100",  "000000000110011011",  "000000000110011010",  "000000000110011001",  "000000000110011000",  "000000000110010111",  "000000000110010110",  "000000000110010100",  "000000000110010011",  "000000000110010010",  "000000000110010001",  "000000000110010000",  "000000000110001111",  "000000000110001110",  "000000000110001100",  "000000000110001011",  "000000000110001010",  "000000000110001001",  "000000000110001000",  "000000000110000111",  "000000000110000101",  "000000000110000100",  "000000000110000011",  "000000000110000010",  "000000000110000001",  "000000000101111111",  "000000000101111110",  "000000000101111101",  "000000000101111100",  "000000000101111011",  "000000000101111001",  "000000000101111000",  "000000000101110111",  "000000000101110110",  "000000000101110100",  "000000000101110011",  "000000000101110010",  "000000000101110001",  "000000000101101111",  "000000000101101110",  "000000000101101101",  "000000000101101100",  "000000000101101010",  "000000000101101001",  "000000000101101000",  "000000000101100110",  "000000000101100101",  "000000000101100100",  "000000000101100011",  "000000000101100001",  "000000000101100000",  "000000000101011111",  "000000000101011101",  "000000000101011100",  "000000000101011011",  "000000000101011001",  "000000000101011000",  "000000000101010111",  "000000000101010101",  "000000000101010100",  "000000000101010011",  "000000000101010001",  "000000000101010000",  "000000000101001111",  "000000000101001101",  "000000000101001100",  "000000000101001011",  "000000000101001001",  "000000000101001000",  "000000000101000110",  "000000000101000101",  "000000000101000100",  "000000000101000010",  "000000000101000001",  "000000000101000000",  "000000000100111110",  "000000000100111101",  "000000000100111011",  "000000000100111010",  "000000000100111001",  "000000000100110111",  "000000000100110110",  "000000000100110100",  "000000000100110011",  "000000000100110001",  "000000000100110000",  "000000000100101111",  "000000000100101101",  "000000000100101100",  "000000000100101010",  "000000000100101001",  "000000000100100111",  "000000000100100110",  "000000000100100100",  "000000000100100011",  "000000000100100001",  "000000000100100000",  "000000000100011110",  "000000000100011101",  "000000000100011100",  "000000000100011010",  "000000000100011001",  "000000000100010111",  "000000000100010110",  "000000000100010100",  "000000000100010011",  "000000000100010001",  "000000000100010000",  "000000000100001110",  "000000000100001101",  "000000000100001011",  "000000000100001001",  "000000000100001000",  "000000000100000110",  "000000000100000101",  "000000000100000011",  "000000000100000010",  "000000000100000000",  "000000000011111111",  "000000000011111101",  "000000000011111100",  "000000000011111010",  "000000000011111001",  "000000000011110111",  "000000000011110101",  "000000000011110100",  "000000000011110010",  "000000000011110001",  "000000000011101111",  "000000000011101110",  "000000000011101100",  "000000000011101010",  "000000000011101001",  "000000000011100111",  "000000000011100110",  "000000000011100100",  "000000000011100010",  "000000000011100001",  "000000000011011111",  "000000000011011110",  "000000000011011100",  "000000000011011010",  "000000000011011001",  "000000000011010111",  "000000000011010110",  "000000000011010100",  "000000000011010010",  "000000000011010001",  "000000000011001111",  "000000000011001101",  "000000000011001100",  "000000000011001010",  "000000000011001000",  "000000000011000111",  "000000000011000101",  "000000000011000100",  "000000000011000010",  "000000000011000000",  "000000000010111111",  "000000000010111101",  "000000000010111011",  "000000000010111010",  "000000000010111000",  "000000000010110110",  "000000000010110101",  "000000000010110011",  "000000000010110001",  "000000000010110000",  "000000000010101110",  "000000000010101100",  "000000000010101011",  "000000000010101001",  "000000000010100111",  "000000000010100101",  "000000000010100100",  "000000000010100010",  "000000000010100000",  "000000000010011111",  "000000000010011101",  "000000000010011011",  "000000000010011010",  "000000000010011000",  "000000000010010110",  "000000000010010100",  "000000000010010011",  "000000000010010001",  "000000000010001111",  "000000000010001110",  "000000000010001100",  "000000000010001010",  "000000000010001000",  "000000000010000111",  "000000000010000101",  "000000000010000011",  "000000000010000001",  "000000000010000000",  "000000000001111110",  "000000000001111100",  "000000000001111010",  "000000000001111001",  "000000000001110111",  "000000000001110101",  "000000000001110011",  "000000000001110010",  "000000000001110000",  "000000000001101110",  "000000000001101100",  "000000000001101011",  "000000000001101001",  "000000000001100111",  "000000000001100101",  "000000000001100100",  "000000000001100010",  "000000000001100000",  "000000000001011110",  "000000000001011100",  "000000000001011011",  "000000000001011001",  "000000000001010111",  "000000000001010101",  "000000000001010100",  "000000000001010010",  "000000000001010000",  "000000000001001110",  "000000000001001100",  "000000000001001011",  "000000000001001001",  "000000000001000111",  "000000000001000101",  "000000000001000011",  "000000000001000010",  "000000000001000000",  "000000000000111110",  "000000000000111100",  "000000000000111010",  "000000000000111001",  "000000000000110111",  "000000000000110101",  "000000000000110011",  "000000000000110001",  "000000000000110000",  "000000000000101110",  "000000000000101100",  "000000000000101010",  "000000000000101000",  "000000000000100110",  "000000000000100101",  "000000000000100011",  "000000000000100001",  "000000000000011111",  "000000000000011101",  "000000000000011100",  "000000000000011010",  "000000000000011000",  "000000000000010110",  "000000000000010100",  "000000000000010010",  "000000000000010001",  "000000000000001111",  "000000000000001101",  "000000000000001011",  "000000000000001001",  "000000000000000111",  "000000000000000110",  "000000000000000100",  "000000000000000010"),("000000000000000000",  "111111111111111110",  "111111111111111100",  "111111111111111010",  "111111111111111001",  "111111111111110111",  "111111111111110101",  "111111111111110011",  "111111111111110001",  "111111111111101111",  "111111111111101110",  "111111111111101100",  "111111111111101010",  "111111111111101000",  "111111111111100110",  "111111111111100100",  "111111111111100010",  "111111111111100001",  "111111111111011111",  "111111111111011101",  "111111111111011011",  "111111111111011001",  "111111111111010111",  "111111111111010101",  "111111111111010100",  "111111111111010010",  "111111111111010000",  "111111111111001110",  "111111111111001100",  "111111111111001010",  "111111111111001001",  "111111111111000111",  "111111111111000101",  "111111111111000011",  "111111111111000001",  "111111111110111111",  "111111111110111101",  "111111111110111100",  "111111111110111010",  "111111111110111000",  "111111111110110110",  "111111111110110100",  "111111111110110010",  "111111111110110000",  "111111111110101110",  "111111111110101101",  "111111111110101011",  "111111111110101001",  "111111111110100111",  "111111111110100101",  "111111111110100011",  "111111111110100001",  "111111111110100000",  "111111111110011110",  "111111111110011100",  "111111111110011010",  "111111111110011000",  "111111111110010110",  "111111111110010100",  "111111111110010011",  "111111111110010001",  "111111111110001111",  "111111111110001101",  "111111111110001011",  "111111111110001001",  "111111111110000111",  "111111111110000110",  "111111111110000100",  "111111111110000010",  "111111111110000000",  "111111111101111110",  "111111111101111100",  "111111111101111011",  "111111111101111001",  "111111111101110111",  "111111111101110101",  "111111111101110011",  "111111111101110001",  "111111111101101111",  "111111111101101110",  "111111111101101100",  "111111111101101010",  "111111111101101000",  "111111111101100110",  "111111111101100100",  "111111111101100010",  "111111111101100001",  "111111111101011111",  "111111111101011101",  "111111111101011011",  "111111111101011001",  "111111111101010111",  "111111111101010110",  "111111111101010100",  "111111111101010010",  "111111111101010000",  "111111111101001110",  "111111111101001100",  "111111111101001011",  "111111111101001001",  "111111111101000111",  "111111111101000101",  "111111111101000011",  "111111111101000001",  "111111111101000000",  "111111111100111110",  "111111111100111100",  "111111111100111010",  "111111111100111000",  "111111111100110110",  "111111111100110101",  "111111111100110011",  "111111111100110001",  "111111111100101111",  "111111111100101101",  "111111111100101100",  "111111111100101010",  "111111111100101000",  "111111111100100110",  "111111111100100100",  "111111111100100010",  "111111111100100001",  "111111111100011111",  "111111111100011101",  "111111111100011011",  "111111111100011001",  "111111111100011000",  "111111111100010110",  "111111111100010100",  "111111111100010010",  "111111111100010000",  "111111111100001111",  "111111111100001101",  "111111111100001011",  "111111111100001001",  "111111111100000111",  "111111111100000110",  "111111111100000100",  "111111111100000010",  "111111111100000000",  "111111111011111111",  "111111111011111101",  "111111111011111011",  "111111111011111001",  "111111111011110111",  "111111111011110110",  "111111111011110100",  "111111111011110010",  "111111111011110000",  "111111111011101111",  "111111111011101101",  "111111111011101011",  "111111111011101001",  "111111111011101000",  "111111111011100110",  "111111111011100100",  "111111111011100010",  "111111111011100001",  "111111111011011111",  "111111111011011101",  "111111111011011011",  "111111111011011010",  "111111111011011000",  "111111111011010110",  "111111111011010100",  "111111111011010011",  "111111111011010001",  "111111111011001111",  "111111111011001101",  "111111111011001100",  "111111111011001010",  "111111111011001000",  "111111111011000111",  "111111111011000101",  "111111111011000011",  "111111111011000001",  "111111111011000000",  "111111111010111110",  "111111111010111100",  "111111111010111011",  "111111111010111001",  "111111111010110111",  "111111111010110101",  "111111111010110100",  "111111111010110010",  "111111111010110000",  "111111111010101111",  "111111111010101101",  "111111111010101011",  "111111111010101010",  "111111111010101000",  "111111111010100110",  "111111111010100101",  "111111111010100011",  "111111111010100001",  "111111111010100000",  "111111111010011110",  "111111111010011100",  "111111111010011011",  "111111111010011001",  "111111111010010111",  "111111111010010110",  "111111111010010100",  "111111111010010010",  "111111111010010001",  "111111111010001111",  "111111111010001110",  "111111111010001100",  "111111111010001010",  "111111111010001001",  "111111111010000111",  "111111111010000101",  "111111111010000100",  "111111111010000010",  "111111111010000001",  "111111111001111111",  "111111111001111101",  "111111111001111100",  "111111111001111010",  "111111111001111001",  "111111111001110111",  "111111111001110101",  "111111111001110100",  "111111111001110010",  "111111111001110001",  "111111111001101111",  "111111111001101101",  "111111111001101100",  "111111111001101010",  "111111111001101001",  "111111111001100111",  "111111111001100110",  "111111111001100100",  "111111111001100011",  "111111111001100001",  "111111111001011111",  "111111111001011110",  "111111111001011100",  "111111111001011011",  "111111111001011001",  "111111111001011000",  "111111111001010110",  "111111111001010101",  "111111111001010011",  "111111111001010010",  "111111111001010000",  "111111111001001111",  "111111111001001101",  "111111111001001100",  "111111111001001010",  "111111111001001001",  "111111111001000111",  "111111111001000110",  "111111111001000100",  "111111111001000011",  "111111111001000001",  "111111111001000000",  "111111111000111110",  "111111111000111101",  "111111111000111011",  "111111111000111010",  "111111111000111000",  "111111111000110111",  "111111111000110110",  "111111111000110100",  "111111111000110011",  "111111111000110001",  "111111111000110000",  "111111111000101110",  "111111111000101101",  "111111111000101100",  "111111111000101010",  "111111111000101001",  "111111111000100111",  "111111111000100110",  "111111111000100100",  "111111111000100011",  "111111111000100010",  "111111111000100000",  "111111111000011111",  "111111111000011110",  "111111111000011100",  "111111111000011011",  "111111111000011001",  "111111111000011000",  "111111111000010111",  "111111111000010101",  "111111111000010100",  "111111111000010011",  "111111111000010001",  "111111111000010000",  "111111111000001111",  "111111111000001101",  "111111111000001100",  "111111111000001011",  "111111111000001001",  "111111111000001000",  "111111111000000111",  "111111111000000101",  "111111111000000100",  "111111111000000011",  "111111111000000001",  "111111111000000000",  "111111110111111111",  "111111110111111110",  "111111110111111100",  "111111110111111011",  "111111110111111010",  "111111110111111000",  "111111110111110111",  "111111110111110110",  "111111110111110101",  "111111110111110011",  "111111110111110010",  "111111110111110001",  "111111110111110000",  "111111110111101111",  "111111110111101101",  "111111110111101100",  "111111110111101011",  "111111110111101010",  "111111110111101000",  "111111110111100111",  "111111110111100110",  "111111110111100101",  "111111110111100100",  "111111110111100010",  "111111110111100001",  "111111110111100000",  "111111110111011111",  "111111110111011110",  "111111110111011101",  "111111110111011011",  "111111110111011010",  "111111110111011001",  "111111110111011000",  "111111110111010111",  "111111110111010110",  "111111110111010101",  "111111110111010011",  "111111110111010010",  "111111110111010001",  "111111110111010000",  "111111110111001111",  "111111110111001110",  "111111110111001101",  "111111110111001100",  "111111110111001011",  "111111110111001010",  "111111110111001001",  "111111110111000111",  "111111110111000110",  "111111110111000101",  "111111110111000100",  "111111110111000011",  "111111110111000010",  "111111110111000001",  "111111110111000000",  "111111110110111111",  "111111110110111110",  "111111110110111101",  "111111110110111100",  "111111110110111011",  "111111110110111010",  "111111110110111001",  "111111110110111000",  "111111110110110111",  "111111110110110110",  "111111110110110101",  "111111110110110100",  "111111110110110011",  "111111110110110010",  "111111110110110001",  "111111110110110000",  "111111110110101111",  "111111110110101110",  "111111110110101101",  "111111110110101100",  "111111110110101100",  "111111110110101011",  "111111110110101010",  "111111110110101001",  "111111110110101000",  "111111110110100111",  "111111110110100110",  "111111110110100101",  "111111110110100100",  "111111110110100011",  "111111110110100011",  "111111110110100010",  "111111110110100001",  "111111110110100000",  "111111110110011111",  "111111110110011110",  "111111110110011101",  "111111110110011101",  "111111110110011100",  "111111110110011011",  "111111110110011010",  "111111110110011001",  "111111110110011000",  "111111110110011000",  "111111110110010111",  "111111110110010110",  "111111110110010101",  "111111110110010101",  "111111110110010100",  "111111110110010011",  "111111110110010010",  "111111110110010001",  "111111110110010001",  "111111110110010000",  "111111110110001111",  "111111110110001110",  "111111110110001110",  "111111110110001101",  "111111110110001100",  "111111110110001100",  "111111110110001011",  "111111110110001010",  "111111110110001001",  "111111110110001001",  "111111110110001000",  "111111110110000111",  "111111110110000111",  "111111110110000110",  "111111110110000101",  "111111110110000101",  "111111110110000100",  "111111110110000011",  "111111110110000011",  "111111110110000010",  "111111110110000010",  "111111110110000001",  "111111110110000000",  "111111110110000000",  "111111110101111111",  "111111110101111110",  "111111110101111110",  "111111110101111101",  "111111110101111101",  "111111110101111100",  "111111110101111100",  "111111110101111011",  "111111110101111010",  "111111110101111010",  "111111110101111001",  "111111110101111001",  "111111110101111000",  "111111110101111000",  "111111110101110111",  "111111110101110111",  "111111110101110110",  "111111110101110110",  "111111110101110101",  "111111110101110101",  "111111110101110100",  "111111110101110100",  "111111110101110011",  "111111110101110011",  "111111110101110010",  "111111110101110010",  "111111110101110001",  "111111110101110001",  "111111110101110000",  "111111110101110000",  "111111110101110000",  "111111110101101111",  "111111110101101111",  "111111110101101110",  "111111110101101110",  "111111110101101110",  "111111110101101101",  "111111110101101101",  "111111110101101100",  "111111110101101100",  "111111110101101100",  "111111110101101011",  "111111110101101011",  "111111110101101011",  "111111110101101010",  "111111110101101010",  "111111110101101010",  "111111110101101001",  "111111110101101001",  "111111110101101001",  "111111110101101000",  "111111110101101000",  "111111110101101000",  "111111110101100111",  "111111110101100111",  "111111110101100111",  "111111110101100111",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100111",  "111111110101100111",  "111111110101100111",  "111111110101101000",  "111111110101101000",  "111111110101101000",  "111111110101101000",  "111111110101101001",  "111111110101101001",  "111111110101101001",  "111111110101101010",  "111111110101101010",  "111111110101101010",  "111111110101101011",  "111111110101101011",  "111111110101101011",  "111111110101101100",  "111111110101101100",  "111111110101101101",  "111111110101101101",  "111111110101101101",  "111111110101101110",  "111111110101101110",  "111111110101101111",  "111111110101101111",  "111111110101101111",  "111111110101110000",  "111111110101110000",  "111111110101110001",  "111111110101110001",  "111111110101110010",  "111111110101110010",  "111111110101110011",  "111111110101110011",  "111111110101110100",  "111111110101110100",  "111111110101110101",  "111111110101110101",  "111111110101110110",  "111111110101110110",  "111111110101110111",  "111111110101110111",  "111111110101111000",  "111111110101111000",  "111111110101111001",  "111111110101111001",  "111111110101111010",  "111111110101111011",  "111111110101111011",  "111111110101111100",  "111111110101111100",  "111111110101111101",  "111111110101111101",  "111111110101111110",  "111111110101111111",  "111111110101111111",  "111111110110000000",  "111111110110000001",  "111111110110000001",  "111111110110000010",  "111111110110000011",  "111111110110000011",  "111111110110000100",  "111111110110000101",  "111111110110000101",  "111111110110000110",  "111111110110000111",  "111111110110000111",  "111111110110001000",  "111111110110001001",  "111111110110001001",  "111111110110001010",  "111111110110001011",  "111111110110001100",  "111111110110001100",  "111111110110001101",  "111111110110001110",  "111111110110001111",  "111111110110001111",  "111111110110010000",  "111111110110010001",  "111111110110010010",  "111111110110010010",  "111111110110010011",  "111111110110010100",  "111111110110010101",  "111111110110010110",  "111111110110010110",  "111111110110010111",  "111111110110011000",  "111111110110011001",  "111111110110011010",  "111111110110011011",  "111111110110011100",  "111111110110011100",  "111111110110011101",  "111111110110011110",  "111111110110011111",  "111111110110100000",  "111111110110100001",  "111111110110100010",  "111111110110100011",  "111111110110100100",  "111111110110100100",  "111111110110100101",  "111111110110100110",  "111111110110100111",  "111111110110101000",  "111111110110101001",  "111111110110101010",  "111111110110101011",  "111111110110101100",  "111111110110101101",  "111111110110101110",  "111111110110101111",  "111111110110110000",  "111111110110110001",  "111111110110110010",  "111111110110110011",  "111111110110110100",  "111111110110110101",  "111111110110110110",  "111111110110110111",  "111111110110111000",  "111111110110111001",  "111111110110111010",  "111111110110111011",  "111111110110111100",  "111111110110111101",  "111111110110111110",  "111111110111000000",  "111111110111000001",  "111111110111000010",  "111111110111000011",  "111111110111000100",  "111111110111000101",  "111111110111000110",  "111111110111000111",  "111111110111001000",  "111111110111001010",  "111111110111001011",  "111111110111001100",  "111111110111001101",  "111111110111001110",  "111111110111001111",  "111111110111010000",  "111111110111010010",  "111111110111010011",  "111111110111010100",  "111111110111010101",  "111111110111010110",  "111111110111011000",  "111111110111011001",  "111111110111011010",  "111111110111011011",  "111111110111011100",  "111111110111011110",  "111111110111011111",  "111111110111100000",  "111111110111100001",  "111111110111100011",  "111111110111100100",  "111111110111100101",  "111111110111100110",  "111111110111101000",  "111111110111101001",  "111111110111101010",  "111111110111101100",  "111111110111101101",  "111111110111101110",  "111111110111110000",  "111111110111110001",  "111111110111110010",  "111111110111110100",  "111111110111110101",  "111111110111110110",  "111111110111111000",  "111111110111111001",  "111111110111111010",  "111111110111111100",  "111111110111111101",  "111111110111111110",  "111111111000000000",  "111111111000000001",  "111111111000000010",  "111111111000000100",  "111111111000000101",  "111111111000000111",  "111111111000001000",  "111111111000001010",  "111111111000001011",  "111111111000001100",  "111111111000001110",  "111111111000001111",  "111111111000010001",  "111111111000010010",  "111111111000010100",  "111111111000010101",  "111111111000010110",  "111111111000011000",  "111111111000011001",  "111111111000011011",  "111111111000011100",  "111111111000011110",  "111111111000011111",  "111111111000100001",  "111111111000100010",  "111111111000100100",  "111111111000100101",  "111111111000100111",  "111111111000101000",  "111111111000101010",  "111111111000101100",  "111111111000101101",  "111111111000101111",  "111111111000110000",  "111111111000110010",  "111111111000110011",  "111111111000110101",  "111111111000110110",  "111111111000111000",  "111111111000111010",  "111111111000111011",  "111111111000111101",  "111111111000111110",  "111111111001000000",  "111111111001000010",  "111111111001000011",  "111111111001000101",  "111111111001000110",  "111111111001001000",  "111111111001001010",  "111111111001001011",  "111111111001001101",  "111111111001001111",  "111111111001010000",  "111111111001010010",  "111111111001010100",  "111111111001010101",  "111111111001010111",  "111111111001011001",  "111111111001011010",  "111111111001011100",  "111111111001011110",  "111111111001011111",  "111111111001100001",  "111111111001100011",  "111111111001100100",  "111111111001100110",  "111111111001101000",  "111111111001101001",  "111111111001101011",  "111111111001101101",  "111111111001101111",  "111111111001110000",  "111111111001110010",  "111111111001110100",  "111111111001110110",  "111111111001110111",  "111111111001111001",  "111111111001111011",  "111111111001111101",  "111111111001111110",  "111111111010000000",  "111111111010000010",  "111111111010000100",  "111111111010000110",  "111111111010000111",  "111111111010001001",  "111111111010001011",  "111111111010001101",  "111111111010001111",  "111111111010010000",  "111111111010010010",  "111111111010010100",  "111111111010010110",  "111111111010011000",  "111111111010011010",  "111111111010011011",  "111111111010011101",  "111111111010011111",  "111111111010100001",  "111111111010100011",  "111111111010100101",  "111111111010100111",  "111111111010101000",  "111111111010101010",  "111111111010101100",  "111111111010101110",  "111111111010110000",  "111111111010110010",  "111111111010110100",  "111111111010110110",  "111111111010111000",  "111111111010111001",  "111111111010111011",  "111111111010111101",  "111111111010111111",  "111111111011000001",  "111111111011000011",  "111111111011000101",  "111111111011000111",  "111111111011001001",  "111111111011001011",  "111111111011001101",  "111111111011001111",  "111111111011010001",  "111111111011010011",  "111111111011010100",  "111111111011010110",  "111111111011011000",  "111111111011011010",  "111111111011011100",  "111111111011011110",  "111111111011100000",  "111111111011100010",  "111111111011100100",  "111111111011100110",  "111111111011101000",  "111111111011101010",  "111111111011101100",  "111111111011101110",  "111111111011110000",  "111111111011110010",  "111111111011110100",  "111111111011110110",  "111111111011111000",  "111111111011111010",  "111111111011111100",  "111111111011111110",  "111111111100000000",  "111111111100000011",  "111111111100000101",  "111111111100000111",  "111111111100001001",  "111111111100001011",  "111111111100001101",  "111111111100001111",  "111111111100010001",  "111111111100010011",  "111111111100010101",  "111111111100010111",  "111111111100011001",  "111111111100011011",  "111111111100011101",  "111111111100011111",  "111111111100100001",  "111111111100100100",  "111111111100100110",  "111111111100101000",  "111111111100101010",  "111111111100101100",  "111111111100101110",  "111111111100110000",  "111111111100110010",  "111111111100110100",  "111111111100110110",  "111111111100111001",  "111111111100111011",  "111111111100111101",  "111111111100111111",  "111111111101000001",  "111111111101000011",  "111111111101000101",  "111111111101000111",  "111111111101001010",  "111111111101001100",  "111111111101001110",  "111111111101010000",  "111111111101010010",  "111111111101010100",  "111111111101010110",  "111111111101011001",  "111111111101011011",  "111111111101011101",  "111111111101011111",  "111111111101100001",  "111111111101100011",  "111111111101100110",  "111111111101101000",  "111111111101101010",  "111111111101101100",  "111111111101101110",  "111111111101110001",  "111111111101110011",  "111111111101110101",  "111111111101110111",  "111111111101111001",  "111111111101111011",  "111111111101111110",  "111111111110000000",  "111111111110000010",  "111111111110000100",  "111111111110000110",  "111111111110001001",  "111111111110001011",  "111111111110001101",  "111111111110001111",  "111111111110010010",  "111111111110010100",  "111111111110010110",  "111111111110011000",  "111111111110011010",  "111111111110011101",  "111111111110011111",  "111111111110100001",  "111111111110100011",  "111111111110100110",  "111111111110101000",  "111111111110101010",  "111111111110101100",  "111111111110101110",  "111111111110110001",  "111111111110110011",  "111111111110110101",  "111111111110110111",  "111111111110111010",  "111111111110111100",  "111111111110111110",  "111111111111000000",  "111111111111000011",  "111111111111000101",  "111111111111000111",  "111111111111001001",  "111111111111001100",  "111111111111001110",  "111111111111010000",  "111111111111010010",  "111111111111010101",  "111111111111010111",  "111111111111011001",  "111111111111011100",  "111111111111011110",  "111111111111100000",  "111111111111100010",  "111111111111100101",  "111111111111100111",  "111111111111101001",  "111111111111101011",  "111111111111101110",  "111111111111110000",  "111111111111110010",  "111111111111110101",  "111111111111110111",  "111111111111111001",  "111111111111111011",  "111111111111111110"),("000000000000000000",  "000000000000000010",  "000000000000000101",  "000000000000000111",  "000000000000001001",  "000000000000001011",  "000000000000001110",  "000000000000010000",  "000000000000010010",  "000000000000010101",  "000000000000010111",  "000000000000011001",  "000000000000011100",  "000000000000011110",  "000000000000100000",  "000000000000100010",  "000000000000100101",  "000000000000100111",  "000000000000101001",  "000000000000101100",  "000000000000101110",  "000000000000110000",  "000000000000110010",  "000000000000110101",  "000000000000110111",  "000000000000111001",  "000000000000111100",  "000000000000111110",  "000000000001000000",  "000000000001000011",  "000000000001000101",  "000000000001000111",  "000000000001001010",  "000000000001001100",  "000000000001001110",  "000000000001010000",  "000000000001010011",  "000000000001010101",  "000000000001010111",  "000000000001011010",  "000000000001011100",  "000000000001011110",  "000000000001100001",  "000000000001100011",  "000000000001100101",  "000000000001101000",  "000000000001101010",  "000000000001101100",  "000000000001101110",  "000000000001110001",  "000000000001110011",  "000000000001110101",  "000000000001111000",  "000000000001111010",  "000000000001111100",  "000000000001111111",  "000000000010000001",  "000000000010000011",  "000000000010000110",  "000000000010001000",  "000000000010001010",  "000000000010001100",  "000000000010001111",  "000000000010010001",  "000000000010010011",  "000000000010010110",  "000000000010011000",  "000000000010011010",  "000000000010011101",  "000000000010011111",  "000000000010100001",  "000000000010100011",  "000000000010100110",  "000000000010101000",  "000000000010101010",  "000000000010101101",  "000000000010101111",  "000000000010110001",  "000000000010110100",  "000000000010110110",  "000000000010111000",  "000000000010111010",  "000000000010111101",  "000000000010111111",  "000000000011000001",  "000000000011000100",  "000000000011000110",  "000000000011001000",  "000000000011001010",  "000000000011001101",  "000000000011001111",  "000000000011010001",  "000000000011010100",  "000000000011010110",  "000000000011011000",  "000000000011011010",  "000000000011011101",  "000000000011011111",  "000000000011100001",  "000000000011100100",  "000000000011100110",  "000000000011101000",  "000000000011101010",  "000000000011101101",  "000000000011101111",  "000000000011110001",  "000000000011110011",  "000000000011110110",  "000000000011111000",  "000000000011111010",  "000000000011111100",  "000000000011111111",  "000000000100000001",  "000000000100000011",  "000000000100000101",  "000000000100001000",  "000000000100001010",  "000000000100001100",  "000000000100001110",  "000000000100010001",  "000000000100010011",  "000000000100010101",  "000000000100010111",  "000000000100011010",  "000000000100011100",  "000000000100011110",  "000000000100100000",  "000000000100100011",  "000000000100100101",  "000000000100100111",  "000000000100101001",  "000000000100101100",  "000000000100101110",  "000000000100110000",  "000000000100110010",  "000000000100110100",  "000000000100110111",  "000000000100111001",  "000000000100111011",  "000000000100111101",  "000000000100111111",  "000000000101000010",  "000000000101000100",  "000000000101000110",  "000000000101001000",  "000000000101001010",  "000000000101001101",  "000000000101001111",  "000000000101010001",  "000000000101010011",  "000000000101010101",  "000000000101011000",  "000000000101011010",  "000000000101011100",  "000000000101011110",  "000000000101100000",  "000000000101100010",  "000000000101100101",  "000000000101100111",  "000000000101101001",  "000000000101101011",  "000000000101101101",  "000000000101101111",  "000000000101110010",  "000000000101110100",  "000000000101110110",  "000000000101111000",  "000000000101111010",  "000000000101111100",  "000000000101111110",  "000000000110000001",  "000000000110000011",  "000000000110000101",  "000000000110000111",  "000000000110001001",  "000000000110001011",  "000000000110001101",  "000000000110001111",  "000000000110010010",  "000000000110010100",  "000000000110010110",  "000000000110011000",  "000000000110011010",  "000000000110011100",  "000000000110011110",  "000000000110100000",  "000000000110100010",  "000000000110100100",  "000000000110100110",  "000000000110101001",  "000000000110101011",  "000000000110101101",  "000000000110101111",  "000000000110110001",  "000000000110110011",  "000000000110110101",  "000000000110110111",  "000000000110111001",  "000000000110111011",  "000000000110111101",  "000000000110111111",  "000000000111000001",  "000000000111000011",  "000000000111000101",  "000000000111000111",  "000000000111001001",  "000000000111001011",  "000000000111001101",  "000000000111001111",  "000000000111010001",  "000000000111010011",  "000000000111010101",  "000000000111010111",  "000000000111011001",  "000000000111011011",  "000000000111011101",  "000000000111011111",  "000000000111100001",  "000000000111100011",  "000000000111100101",  "000000000111100111",  "000000000111101001",  "000000000111101011",  "000000000111101101",  "000000000111101111",  "000000000111110001",  "000000000111110011",  "000000000111110101",  "000000000111110111",  "000000000111111001",  "000000000111111011",  "000000000111111101",  "000000000111111111",  "000000001000000001",  "000000001000000010",  "000000001000000100",  "000000001000000110",  "000000001000001000",  "000000001000001010",  "000000001000001100",  "000000001000001110",  "000000001000010000",  "000000001000010010",  "000000001000010100",  "000000001000010101",  "000000001000010111",  "000000001000011001",  "000000001000011011",  "000000001000011101",  "000000001000011111",  "000000001000100001",  "000000001000100010",  "000000001000100100",  "000000001000100110",  "000000001000101000",  "000000001000101010",  "000000001000101100",  "000000001000101101",  "000000001000101111",  "000000001000110001",  "000000001000110011",  "000000001000110101",  "000000001000110110",  "000000001000111000",  "000000001000111010",  "000000001000111100",  "000000001000111101",  "000000001000111111",  "000000001001000001",  "000000001001000011",  "000000001001000101",  "000000001001000110",  "000000001001001000",  "000000001001001010",  "000000001001001011",  "000000001001001101",  "000000001001001111",  "000000001001010001",  "000000001001010010",  "000000001001010100",  "000000001001010110",  "000000001001011000",  "000000001001011001",  "000000001001011011",  "000000001001011101",  "000000001001011110",  "000000001001100000",  "000000001001100010",  "000000001001100011",  "000000001001100101",  "000000001001100111",  "000000001001101000",  "000000001001101010",  "000000001001101100",  "000000001001101101",  "000000001001101111",  "000000001001110000",  "000000001001110010",  "000000001001110100",  "000000001001110101",  "000000001001110111",  "000000001001111000",  "000000001001111010",  "000000001001111100",  "000000001001111101",  "000000001001111111",  "000000001010000000",  "000000001010000010",  "000000001010000100",  "000000001010000101",  "000000001010000111",  "000000001010001000",  "000000001010001010",  "000000001010001011",  "000000001010001101",  "000000001010001110",  "000000001010010000",  "000000001010010001",  "000000001010010011",  "000000001010010100",  "000000001010010110",  "000000001010010111",  "000000001010011001",  "000000001010011010",  "000000001010011100",  "000000001010011101",  "000000001010011111",  "000000001010100000",  "000000001010100010",  "000000001010100011",  "000000001010100100",  "000000001010100110",  "000000001010100111",  "000000001010101001",  "000000001010101010",  "000000001010101100",  "000000001010101101",  "000000001010101110",  "000000001010110000",  "000000001010110001",  "000000001010110010",  "000000001010110100",  "000000001010110101",  "000000001010110111",  "000000001010111000",  "000000001010111001",  "000000001010111011",  "000000001010111100",  "000000001010111101",  "000000001010111111",  "000000001011000000",  "000000001011000001",  "000000001011000011",  "000000001011000100",  "000000001011000101",  "000000001011000110",  "000000001011001000",  "000000001011001001",  "000000001011001010",  "000000001011001100",  "000000001011001101",  "000000001011001110",  "000000001011001111",  "000000001011010001",  "000000001011010010",  "000000001011010011",  "000000001011010100",  "000000001011010101",  "000000001011010111",  "000000001011011000",  "000000001011011001",  "000000001011011010",  "000000001011011011",  "000000001011011101",  "000000001011011110",  "000000001011011111",  "000000001011100000",  "000000001011100001",  "000000001011100010",  "000000001011100011",  "000000001011100101",  "000000001011100110",  "000000001011100111",  "000000001011101000",  "000000001011101001",  "000000001011101010",  "000000001011101011",  "000000001011101100",  "000000001011101101",  "000000001011101110",  "000000001011101111",  "000000001011110001",  "000000001011110010",  "000000001011110011",  "000000001011110100",  "000000001011110101",  "000000001011110110",  "000000001011110111",  "000000001011111000",  "000000001011111001",  "000000001011111010",  "000000001011111011",  "000000001011111100",  "000000001011111101",  "000000001011111110",  "000000001011111111",  "000000001100000000",  "000000001100000001",  "000000001100000001",  "000000001100000010",  "000000001100000011",  "000000001100000100",  "000000001100000101",  "000000001100000110",  "000000001100000111",  "000000001100001000",  "000000001100001001",  "000000001100001010",  "000000001100001010",  "000000001100001011",  "000000001100001100",  "000000001100001101",  "000000001100001110",  "000000001100001111",  "000000001100010000",  "000000001100010000",  "000000001100010001",  "000000001100010010",  "000000001100010011",  "000000001100010100",  "000000001100010100",  "000000001100010101",  "000000001100010110",  "000000001100010111",  "000000001100010111",  "000000001100011000",  "000000001100011001",  "000000001100011010",  "000000001100011010",  "000000001100011011",  "000000001100011100",  "000000001100011101",  "000000001100011101",  "000000001100011110",  "000000001100011111",  "000000001100011111",  "000000001100100000",  "000000001100100001",  "000000001100100001",  "000000001100100010",  "000000001100100011",  "000000001100100011",  "000000001100100100",  "000000001100100100",  "000000001100100101",  "000000001100100110",  "000000001100100110",  "000000001100100111",  "000000001100100111",  "000000001100101000",  "000000001100101001",  "000000001100101001",  "000000001100101010",  "000000001100101010",  "000000001100101011",  "000000001100101011",  "000000001100101100",  "000000001100101100",  "000000001100101101",  "000000001100101101",  "000000001100101110",  "000000001100101110",  "000000001100101111",  "000000001100101111",  "000000001100110000",  "000000001100110000",  "000000001100110001",  "000000001100110001",  "000000001100110001",  "000000001100110010",  "000000001100110010",  "000000001100110011",  "000000001100110011",  "000000001100110100",  "000000001100110100",  "000000001100110100",  "000000001100110101",  "000000001100110101",  "000000001100110101",  "000000001100110110",  "000000001100110110",  "000000001100110110",  "000000001100110111",  "000000001100110111",  "000000001100110111",  "000000001100111000",  "000000001100111000",  "000000001100111000",  "000000001100111001",  "000000001100111001",  "000000001100111001",  "000000001100111001",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111001",  "000000001100111001",  "000000001100111001",  "000000001100111000",  "000000001100111000",  "000000001100111000",  "000000001100111000",  "000000001100110111",  "000000001100110111",  "000000001100110111",  "000000001100110110",  "000000001100110110",  "000000001100110110",  "000000001100110101",  "000000001100110101",  "000000001100110101",  "000000001100110100",  "000000001100110100",  "000000001100110011",  "000000001100110011",  "000000001100110011",  "000000001100110010",  "000000001100110010",  "000000001100110001",  "000000001100110001",  "000000001100110000",  "000000001100110000",  "000000001100101111",  "000000001100101111",  "000000001100101111",  "000000001100101110",  "000000001100101110",  "000000001100101101",  "000000001100101100",  "000000001100101100",  "000000001100101011",  "000000001100101011",  "000000001100101010",  "000000001100101010",  "000000001100101001",  "000000001100101001",  "000000001100101000",  "000000001100101000",  "000000001100100111",  "000000001100100110",  "000000001100100110",  "000000001100100101",  "000000001100100100",  "000000001100100100",  "000000001100100011",  "000000001100100011",  "000000001100100010",  "000000001100100001",  "000000001100100001",  "000000001100100000",  "000000001100011111",  "000000001100011111",  "000000001100011110",  "000000001100011101",  "000000001100011100",  "000000001100011100",  "000000001100011011",  "000000001100011010",  "000000001100011001",  "000000001100011001",  "000000001100011000",  "000000001100010111",  "000000001100010110",  "000000001100010110",  "000000001100010101",  "000000001100010100",  "000000001100010011",  "000000001100010010",  "000000001100010001",  "000000001100010001",  "000000001100010000",  "000000001100001111",  "000000001100001110",  "000000001100001101",  "000000001100001100",  "000000001100001011",  "000000001100001011",  "000000001100001010",  "000000001100001001",  "000000001100001000",  "000000001100000111",  "000000001100000110",  "000000001100000101",  "000000001100000100",  "000000001100000011",  "000000001100000010",  "000000001100000001",  "000000001100000000",  "000000001011111111",  "000000001011111110",  "000000001011111101",  "000000001011111100",  "000000001011111011",  "000000001011111010",  "000000001011111001",  "000000001011111000",  "000000001011110111",  "000000001011110110",  "000000001011110101",  "000000001011110100",  "000000001011110011",  "000000001011110010",  "000000001011110001",  "000000001011110000",  "000000001011101111",  "000000001011101101",  "000000001011101100",  "000000001011101011",  "000000001011101010",  "000000001011101001",  "000000001011101000",  "000000001011100111",  "000000001011100101",  "000000001011100100",  "000000001011100011",  "000000001011100010",  "000000001011100001",  "000000001011100000",  "000000001011011110",  "000000001011011101",  "000000001011011100",  "000000001011011011",  "000000001011011001",  "000000001011011000",  "000000001011010111",  "000000001011010110",  "000000001011010100",  "000000001011010011",  "000000001011010010",  "000000001011010001",  "000000001011001111",  "000000001011001110",  "000000001011001101",  "000000001011001011",  "000000001011001010",  "000000001011001001",  "000000001011000111",  "000000001011000110",  "000000001011000101",  "000000001011000011",  "000000001011000010",  "000000001011000001",  "000000001010111111",  "000000001010111110",  "000000001010111100",  "000000001010111011",  "000000001010111010",  "000000001010111000",  "000000001010110111",  "000000001010110101",  "000000001010110100",  "000000001010110010",  "000000001010110001",  "000000001010101111",  "000000001010101110",  "000000001010101100",  "000000001010101011",  "000000001010101010",  "000000001010101000",  "000000001010100110",  "000000001010100101",  "000000001010100011",  "000000001010100010",  "000000001010100000",  "000000001010011111",  "000000001010011101",  "000000001010011100",  "000000001010011010",  "000000001010011001",  "000000001010010111",  "000000001010010101",  "000000001010010100",  "000000001010010010",  "000000001010010001",  "000000001010001111",  "000000001010001101",  "000000001010001100",  "000000001010001010",  "000000001010001001",  "000000001010000111",  "000000001010000101",  "000000001010000100",  "000000001010000010",  "000000001010000000",  "000000001001111111",  "000000001001111101",  "000000001001111011",  "000000001001111010",  "000000001001111000",  "000000001001110110",  "000000001001110100",  "000000001001110011",  "000000001001110001",  "000000001001101111",  "000000001001101101",  "000000001001101100",  "000000001001101010",  "000000001001101000",  "000000001001100110",  "000000001001100101",  "000000001001100011",  "000000001001100001",  "000000001001011111",  "000000001001011101",  "000000001001011100",  "000000001001011010",  "000000001001011000",  "000000001001010110",  "000000001001010100",  "000000001001010011",  "000000001001010001",  "000000001001001111",  "000000001001001101",  "000000001001001011",  "000000001001001001",  "000000001001000111",  "000000001001000101",  "000000001001000100",  "000000001001000010",  "000000001001000000",  "000000001000111110",  "000000001000111100",  "000000001000111010",  "000000001000111000",  "000000001000110110",  "000000001000110100",  "000000001000110010",  "000000001000110000",  "000000001000101110",  "000000001000101100",  "000000001000101010",  "000000001000101000",  "000000001000100110",  "000000001000100100",  "000000001000100010",  "000000001000100000",  "000000001000011110",  "000000001000011100",  "000000001000011010",  "000000001000011000",  "000000001000010110",  "000000001000010100",  "000000001000010010",  "000000001000010000",  "000000001000001110",  "000000001000001100",  "000000001000001010",  "000000001000001000",  "000000001000000110",  "000000001000000100",  "000000001000000010",  "000000001000000000",  "000000000111111110",  "000000000111111011",  "000000000111111001",  "000000000111110111",  "000000000111110101",  "000000000111110011",  "000000000111110001",  "000000000111101111",  "000000000111101101",  "000000000111101010",  "000000000111101000",  "000000000111100110",  "000000000111100100",  "000000000111100010",  "000000000111100000",  "000000000111011101",  "000000000111011011",  "000000000111011001",  "000000000111010111",  "000000000111010101",  "000000000111010010",  "000000000111010000",  "000000000111001110",  "000000000111001100",  "000000000111001001",  "000000000111000111",  "000000000111000101",  "000000000111000011",  "000000000111000000",  "000000000110111110",  "000000000110111100",  "000000000110111010",  "000000000110110111",  "000000000110110101",  "000000000110110011",  "000000000110110001",  "000000000110101110",  "000000000110101100",  "000000000110101010",  "000000000110100111",  "000000000110100101",  "000000000110100011",  "000000000110100000",  "000000000110011110",  "000000000110011100",  "000000000110011001",  "000000000110010111",  "000000000110010101",  "000000000110010010",  "000000000110010000",  "000000000110001110",  "000000000110001011",  "000000000110001001",  "000000000110000111",  "000000000110000100",  "000000000110000010",  "000000000101111111",  "000000000101111101",  "000000000101111011",  "000000000101111000",  "000000000101110110",  "000000000101110011",  "000000000101110001",  "000000000101101111",  "000000000101101100",  "000000000101101010",  "000000000101100111",  "000000000101100101",  "000000000101100010",  "000000000101100000",  "000000000101011110",  "000000000101011011",  "000000000101011001",  "000000000101010110",  "000000000101010100",  "000000000101010001",  "000000000101001111",  "000000000101001100",  "000000000101001010",  "000000000101000111",  "000000000101000101",  "000000000101000010",  "000000000101000000",  "000000000100111101",  "000000000100111011",  "000000000100111000",  "000000000100110110",  "000000000100110011",  "000000000100110001",  "000000000100101110",  "000000000100101100",  "000000000100101001",  "000000000100100111",  "000000000100100100",  "000000000100100001",  "000000000100011111",  "000000000100011100",  "000000000100011010",  "000000000100010111",  "000000000100010101",  "000000000100010010",  "000000000100010000",  "000000000100001101",  "000000000100001010",  "000000000100001000",  "000000000100000101",  "000000000100000011",  "000000000100000000",  "000000000011111101",  "000000000011111011",  "000000000011111000",  "000000000011110110",  "000000000011110011",  "000000000011110000",  "000000000011101110",  "000000000011101011",  "000000000011101000",  "000000000011100110",  "000000000011100011",  "000000000011100001",  "000000000011011110",  "000000000011011011",  "000000000011011001",  "000000000011010110",  "000000000011010011",  "000000000011010001",  "000000000011001110",  "000000000011001011",  "000000000011001001",  "000000000011000110",  "000000000011000011",  "000000000011000001",  "000000000010111110",  "000000000010111011",  "000000000010111001",  "000000000010110110",  "000000000010110011",  "000000000010110001",  "000000000010101110",  "000000000010101011",  "000000000010101001",  "000000000010100110",  "000000000010100011",  "000000000010100000",  "000000000010011110",  "000000000010011011",  "000000000010011000",  "000000000010010110",  "000000000010010011",  "000000000010010000",  "000000000010001101",  "000000000010001011",  "000000000010001000",  "000000000010000101",  "000000000010000011",  "000000000010000000",  "000000000001111101",  "000000000001111010",  "000000000001111000",  "000000000001110101",  "000000000001110010",  "000000000001101111",  "000000000001101101",  "000000000001101010",  "000000000001100111",  "000000000001100100",  "000000000001100010",  "000000000001011111",  "000000000001011100",  "000000000001011001",  "000000000001010111",  "000000000001010100",  "000000000001010001",  "000000000001001110",  "000000000001001011",  "000000000001001001",  "000000000001000110",  "000000000001000011",  "000000000001000000",  "000000000000111110",  "000000000000111011",  "000000000000111000",  "000000000000110101",  "000000000000110010",  "000000000000110000",  "000000000000101101",  "000000000000101010",  "000000000000100111",  "000000000000100100",  "000000000000100010",  "000000000000011111",  "000000000000011100",  "000000000000011001",  "000000000000010110",  "000000000000010100",  "000000000000010001",  "000000000000001110",  "000000000000001011",  "000000000000001000",  "000000000000000110",  "000000000000000011"),("000000000000000000",  "111111111111111101",  "111111111111111010",  "111111111111111000",  "111111111111110101",  "111111111111110010",  "111111111111101111",  "111111111111101100",  "111111111111101001",  "111111111111100111",  "111111111111100100",  "111111111111100001",  "111111111111011110",  "111111111111011011",  "111111111111011001",  "111111111111010110",  "111111111111010011",  "111111111111010000",  "111111111111001101",  "111111111111001010",  "111111111111001000",  "111111111111000101",  "111111111111000010",  "111111111110111111",  "111111111110111100",  "111111111110111001",  "111111111110110111",  "111111111110110100",  "111111111110110001",  "111111111110101110",  "111111111110101011",  "111111111110101000",  "111111111110100110",  "111111111110100011",  "111111111110100000",  "111111111110011101",  "111111111110011010",  "111111111110010111",  "111111111110010101",  "111111111110010010",  "111111111110001111",  "111111111110001100",  "111111111110001001",  "111111111110000110",  "111111111110000100",  "111111111110000001",  "111111111101111110",  "111111111101111011",  "111111111101111000",  "111111111101110101",  "111111111101110010",  "111111111101110000",  "111111111101101101",  "111111111101101010",  "111111111101100111",  "111111111101100100",  "111111111101100001",  "111111111101011111",  "111111111101011100",  "111111111101011001",  "111111111101010110",  "111111111101010011",  "111111111101010000",  "111111111101001110",  "111111111101001011",  "111111111101001000",  "111111111101000101",  "111111111101000010",  "111111111100111111",  "111111111100111101",  "111111111100111010",  "111111111100110111",  "111111111100110100",  "111111111100110001",  "111111111100101111",  "111111111100101100",  "111111111100101001",  "111111111100100110",  "111111111100100011",  "111111111100100000",  "111111111100011110",  "111111111100011011",  "111111111100011000",  "111111111100010101",  "111111111100010010",  "111111111100010000",  "111111111100001101",  "111111111100001010",  "111111111100000111",  "111111111100000100",  "111111111100000001",  "111111111011111111",  "111111111011111100",  "111111111011111001",  "111111111011110110",  "111111111011110011",  "111111111011110001",  "111111111011101110",  "111111111011101011",  "111111111011101000",  "111111111011100110",  "111111111011100011",  "111111111011100000",  "111111111011011101",  "111111111011011010",  "111111111011011000",  "111111111011010101",  "111111111011010010",  "111111111011001111",  "111111111011001100",  "111111111011001010",  "111111111011000111",  "111111111011000100",  "111111111011000001",  "111111111010111111",  "111111111010111100",  "111111111010111001",  "111111111010110110",  "111111111010110100",  "111111111010110001",  "111111111010101110",  "111111111010101011",  "111111111010101001",  "111111111010100110",  "111111111010100011",  "111111111010100000",  "111111111010011110",  "111111111010011011",  "111111111010011000",  "111111111010010101",  "111111111010010011",  "111111111010010000",  "111111111010001101",  "111111111010001010",  "111111111010001000",  "111111111010000101",  "111111111010000010",  "111111111010000000",  "111111111001111101",  "111111111001111010",  "111111111001110111",  "111111111001110101",  "111111111001110010",  "111111111001101111",  "111111111001101101",  "111111111001101010",  "111111111001100111",  "111111111001100101",  "111111111001100010",  "111111111001011111",  "111111111001011100",  "111111111001011010",  "111111111001010111",  "111111111001010100",  "111111111001010010",  "111111111001001111",  "111111111001001100",  "111111111001001010",  "111111111001000111",  "111111111001000100",  "111111111001000010",  "111111111000111111",  "111111111000111101",  "111111111000111010",  "111111111000110111",  "111111111000110101",  "111111111000110010",  "111111111000101111",  "111111111000101101",  "111111111000101010",  "111111111000100111",  "111111111000100101",  "111111111000100010",  "111111111000100000",  "111111111000011101",  "111111111000011010",  "111111111000011000",  "111111111000010101",  "111111111000010011",  "111111111000010000",  "111111111000001101",  "111111111000001011",  "111111111000001000",  "111111111000000110",  "111111111000000011",  "111111111000000001",  "111111110111111110",  "111111110111111100",  "111111110111111001",  "111111110111110110",  "111111110111110100",  "111111110111110001",  "111111110111101111",  "111111110111101100",  "111111110111101010",  "111111110111100111",  "111111110111100101",  "111111110111100010",  "111111110111100000",  "111111110111011101",  "111111110111011011",  "111111110111011000",  "111111110111010110",  "111111110111010011",  "111111110111010001",  "111111110111001110",  "111111110111001100",  "111111110111001001",  "111111110111000111",  "111111110111000100",  "111111110111000010",  "111111110110111111",  "111111110110111101",  "111111110110111011",  "111111110110111000",  "111111110110110110",  "111111110110110011",  "111111110110110001",  "111111110110101110",  "111111110110101100",  "111111110110101010",  "111111110110100111",  "111111110110100101",  "111111110110100010",  "111111110110100000",  "111111110110011110",  "111111110110011011",  "111111110110011001",  "111111110110010110",  "111111110110010100",  "111111110110010010",  "111111110110001111",  "111111110110001101",  "111111110110001011",  "111111110110001000",  "111111110110000110",  "111111110110000100",  "111111110110000001",  "111111110101111111",  "111111110101111101",  "111111110101111010",  "111111110101111000",  "111111110101110110",  "111111110101110011",  "111111110101110001",  "111111110101101111",  "111111110101101100",  "111111110101101010",  "111111110101101000",  "111111110101100110",  "111111110101100011",  "111111110101100001",  "111111110101011111",  "111111110101011101",  "111111110101011010",  "111111110101011000",  "111111110101010110",  "111111110101010100",  "111111110101010001",  "111111110101001111",  "111111110101001101",  "111111110101001011",  "111111110101001001",  "111111110101000110",  "111111110101000100",  "111111110101000010",  "111111110101000000",  "111111110100111110",  "111111110100111100",  "111111110100111001",  "111111110100110111",  "111111110100110101",  "111111110100110011",  "111111110100110001",  "111111110100101111",  "111111110100101101",  "111111110100101011",  "111111110100101000",  "111111110100100110",  "111111110100100100",  "111111110100100010",  "111111110100100000",  "111111110100011110",  "111111110100011100",  "111111110100011010",  "111111110100011000",  "111111110100010110",  "111111110100010100",  "111111110100010010",  "111111110100010000",  "111111110100001110",  "111111110100001100",  "111111110100001010",  "111111110100001000",  "111111110100000110",  "111111110100000100",  "111111110100000010",  "111111110100000000",  "111111110011111110",  "111111110011111100",  "111111110011111010",  "111111110011111000",  "111111110011110110",  "111111110011110100",  "111111110011110010",  "111111110011110000",  "111111110011101110",  "111111110011101100",  "111111110011101010",  "111111110011101000",  "111111110011100110",  "111111110011100101",  "111111110011100011",  "111111110011100001",  "111111110011011111",  "111111110011011101",  "111111110011011011",  "111111110011011001",  "111111110011011000",  "111111110011010110",  "111111110011010100",  "111111110011010010",  "111111110011010000",  "111111110011001110",  "111111110011001101",  "111111110011001011",  "111111110011001001",  "111111110011000111",  "111111110011000101",  "111111110011000100",  "111111110011000010",  "111111110011000000",  "111111110010111110",  "111111110010111101",  "111111110010111011",  "111111110010111001",  "111111110010111000",  "111111110010110110",  "111111110010110100",  "111111110010110010",  "111111110010110001",  "111111110010101111",  "111111110010101101",  "111111110010101100",  "111111110010101010",  "111111110010101000",  "111111110010100111",  "111111110010100101",  "111111110010100100",  "111111110010100010",  "111111110010100000",  "111111110010011111",  "111111110010011101",  "111111110010011100",  "111111110010011010",  "111111110010011000",  "111111110010010111",  "111111110010010101",  "111111110010010100",  "111111110010010010",  "111111110010010001",  "111111110010001111",  "111111110010001110",  "111111110010001100",  "111111110010001011",  "111111110010001001",  "111111110010001000",  "111111110010000110",  "111111110010000101",  "111111110010000011",  "111111110010000010",  "111111110010000000",  "111111110001111111",  "111111110001111101",  "111111110001111100",  "111111110001111011",  "111111110001111001",  "111111110001111000",  "111111110001110110",  "111111110001110101",  "111111110001110100",  "111111110001110010",  "111111110001110001",  "111111110001110000",  "111111110001101110",  "111111110001101101",  "111111110001101100",  "111111110001101010",  "111111110001101001",  "111111110001101000",  "111111110001100110",  "111111110001100101",  "111111110001100100",  "111111110001100010",  "111111110001100001",  "111111110001100000",  "111111110001011111",  "111111110001011101",  "111111110001011100",  "111111110001011011",  "111111110001011010",  "111111110001011001",  "111111110001010111",  "111111110001010110",  "111111110001010101",  "111111110001010100",  "111111110001010011",  "111111110001010010",  "111111110001010000",  "111111110001001111",  "111111110001001110",  "111111110001001101",  "111111110001001100",  "111111110001001011",  "111111110001001010",  "111111110001001001",  "111111110001001000",  "111111110001000111",  "111111110001000101",  "111111110001000100",  "111111110001000011",  "111111110001000010",  "111111110001000001",  "111111110001000000",  "111111110000111111",  "111111110000111110",  "111111110000111101",  "111111110000111100",  "111111110000111011",  "111111110000111010",  "111111110000111001",  "111111110000111000",  "111111110000111000",  "111111110000110111",  "111111110000110110",  "111111110000110101",  "111111110000110100",  "111111110000110011",  "111111110000110010",  "111111110000110001",  "111111110000110000",  "111111110000101111",  "111111110000101111",  "111111110000101110",  "111111110000101101",  "111111110000101100",  "111111110000101011",  "111111110000101011",  "111111110000101010",  "111111110000101001",  "111111110000101000",  "111111110000100111",  "111111110000100111",  "111111110000100110",  "111111110000100101",  "111111110000100100",  "111111110000100100",  "111111110000100011",  "111111110000100010",  "111111110000100010",  "111111110000100001",  "111111110000100000",  "111111110000100000",  "111111110000011111",  "111111110000011110",  "111111110000011110",  "111111110000011101",  "111111110000011100",  "111111110000011100",  "111111110000011011",  "111111110000011011",  "111111110000011010",  "111111110000011001",  "111111110000011001",  "111111110000011000",  "111111110000011000",  "111111110000010111",  "111111110000010111",  "111111110000010110",  "111111110000010110",  "111111110000010101",  "111111110000010101",  "111111110000010100",  "111111110000010100",  "111111110000010011",  "111111110000010011",  "111111110000010010",  "111111110000010010",  "111111110000010001",  "111111110000010001",  "111111110000010001",  "111111110000010000",  "111111110000010000",  "111111110000001111",  "111111110000001111",  "111111110000001111",  "111111110000001110",  "111111110000001110",  "111111110000001110",  "111111110000001101",  "111111110000001101",  "111111110000001101",  "111111110000001100",  "111111110000001100",  "111111110000001100",  "111111110000001100",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001100",  "111111110000001100",  "111111110000001100",  "111111110000001101",  "111111110000001101",  "111111110000001101",  "111111110000001110",  "111111110000001110",  "111111110000001110",  "111111110000001111",  "111111110000001111",  "111111110000001111",  "111111110000010000",  "111111110000010000",  "111111110000010001",  "111111110000010001",  "111111110000010001",  "111111110000010010",  "111111110000010010",  "111111110000010011",  "111111110000010011",  "111111110000010100",  "111111110000010100",  "111111110000010101",  "111111110000010101",  "111111110000010110",  "111111110000010110",  "111111110000010111",  "111111110000010111",  "111111110000011000",  "111111110000011000",  "111111110000011001",  "111111110000011001",  "111111110000011010",  "111111110000011011",  "111111110000011011",  "111111110000011100",  "111111110000011101",  "111111110000011101",  "111111110000011110",  "111111110000011110",  "111111110000011111",  "111111110000100000",  "111111110000100000",  "111111110000100001",  "111111110000100010",  "111111110000100011",  "111111110000100011",  "111111110000100100",  "111111110000100101",  "111111110000100110",  "111111110000100110",  "111111110000100111",  "111111110000101000",  "111111110000101001",  "111111110000101001",  "111111110000101010",  "111111110000101011",  "111111110000101100",  "111111110000101101",  "111111110000101110",  "111111110000101110",  "111111110000101111",  "111111110000110000",  "111111110000110001",  "111111110000110010",  "111111110000110011",  "111111110000110100",  "111111110000110101",  "111111110000110110",  "111111110000110111",  "111111110000111000",  "111111110000111001",  "111111110000111001",  "111111110000111010",  "111111110000111011",  "111111110000111100",  "111111110000111101",  "111111110000111111",  "111111110001000000",  "111111110001000001",  "111111110001000010",  "111111110001000011",  "111111110001000100",  "111111110001000101",  "111111110001000110",  "111111110001000111",  "111111110001001000",  "111111110001001001",  "111111110001001010",  "111111110001001011",  "111111110001001101",  "111111110001001110",  "111111110001001111",  "111111110001010000",  "111111110001010001",  "111111110001010010",  "111111110001010100",  "111111110001010101",  "111111110001010110",  "111111110001010111",  "111111110001011001",  "111111110001011010",  "111111110001011011",  "111111110001011100",  "111111110001011110",  "111111110001011111",  "111111110001100000",  "111111110001100001",  "111111110001100011",  "111111110001100100",  "111111110001100101",  "111111110001100111",  "111111110001101000",  "111111110001101010",  "111111110001101011",  "111111110001101100",  "111111110001101110",  "111111110001101111",  "111111110001110000",  "111111110001110010",  "111111110001110011",  "111111110001110101",  "111111110001110110",  "111111110001111000",  "111111110001111001",  "111111110001111011",  "111111110001111100",  "111111110001111101",  "111111110001111111",  "111111110010000000",  "111111110010000010",  "111111110010000100",  "111111110010000101",  "111111110010000111",  "111111110010001000",  "111111110010001010",  "111111110010001011",  "111111110010001101",  "111111110010001110",  "111111110010010000",  "111111110010010010",  "111111110010010011",  "111111110010010101",  "111111110010010110",  "111111110010011000",  "111111110010011010",  "111111110010011011",  "111111110010011101",  "111111110010011111",  "111111110010100000",  "111111110010100010",  "111111110010100100",  "111111110010100110",  "111111110010100111",  "111111110010101001",  "111111110010101011",  "111111110010101100",  "111111110010101110",  "111111110010110000",  "111111110010110010",  "111111110010110100",  "111111110010110101",  "111111110010110111",  "111111110010111001",  "111111110010111011",  "111111110010111101",  "111111110010111110",  "111111110011000000",  "111111110011000010",  "111111110011000100",  "111111110011000110",  "111111110011001000",  "111111110011001010",  "111111110011001011",  "111111110011001101",  "111111110011001111",  "111111110011010001",  "111111110011010011",  "111111110011010101",  "111111110011010111",  "111111110011011001",  "111111110011011011",  "111111110011011101",  "111111110011011111",  "111111110011100001",  "111111110011100011",  "111111110011100101",  "111111110011100111",  "111111110011101001",  "111111110011101011",  "111111110011101101",  "111111110011101111",  "111111110011110001",  "111111110011110011",  "111111110011110101",  "111111110011110111",  "111111110011111001",  "111111110011111011",  "111111110011111101",  "111111110100000000",  "111111110100000010",  "111111110100000100",  "111111110100000110",  "111111110100001000",  "111111110100001010",  "111111110100001100",  "111111110100001110",  "111111110100010001",  "111111110100010011",  "111111110100010101",  "111111110100010111",  "111111110100011001",  "111111110100011100",  "111111110100011110",  "111111110100100000",  "111111110100100010",  "111111110100100101",  "111111110100100111",  "111111110100101001",  "111111110100101011",  "111111110100101110",  "111111110100110000",  "111111110100110010",  "111111110100110100",  "111111110100110111",  "111111110100111001",  "111111110100111011",  "111111110100111110",  "111111110101000000",  "111111110101000010",  "111111110101000101",  "111111110101000111",  "111111110101001001",  "111111110101001100",  "111111110101001110",  "111111110101010001",  "111111110101010011",  "111111110101010101",  "111111110101011000",  "111111110101011010",  "111111110101011101",  "111111110101011111",  "111111110101100001",  "111111110101100100",  "111111110101100110",  "111111110101101001",  "111111110101101011",  "111111110101101110",  "111111110101110000",  "111111110101110011",  "111111110101110101",  "111111110101111000",  "111111110101111010",  "111111110101111101",  "111111110101111111",  "111111110110000010",  "111111110110000100",  "111111110110000111",  "111111110110001001",  "111111110110001100",  "111111110110001111",  "111111110110010001",  "111111110110010100",  "111111110110010110",  "111111110110011001",  "111111110110011100",  "111111110110011110",  "111111110110100001",  "111111110110100011",  "111111110110100110",  "111111110110101001",  "111111110110101011",  "111111110110101110",  "111111110110110001",  "111111110110110011",  "111111110110110110",  "111111110110111001",  "111111110110111011",  "111111110110111110",  "111111110111000001",  "111111110111000011",  "111111110111000110",  "111111110111001001",  "111111110111001011",  "111111110111001110",  "111111110111010001",  "111111110111010100",  "111111110111010110",  "111111110111011001",  "111111110111011100",  "111111110111011111",  "111111110111100001",  "111111110111100100",  "111111110111100111",  "111111110111101010",  "111111110111101101",  "111111110111101111",  "111111110111110010",  "111111110111110101",  "111111110111111000",  "111111110111111011",  "111111110111111101",  "111111111000000000",  "111111111000000011",  "111111111000000110",  "111111111000001001",  "111111111000001100",  "111111111000001111",  "111111111000010001",  "111111111000010100",  "111111111000010111",  "111111111000011010",  "111111111000011101",  "111111111000100000",  "111111111000100011",  "111111111000100110",  "111111111000101001",  "111111111000101100",  "111111111000101110",  "111111111000110001",  "111111111000110100",  "111111111000110111",  "111111111000111010",  "111111111000111101",  "111111111001000000",  "111111111001000011",  "111111111001000110",  "111111111001001001",  "111111111001001100",  "111111111001001111",  "111111111001010010",  "111111111001010101",  "111111111001011000",  "111111111001011011",  "111111111001011110",  "111111111001100001",  "111111111001100100",  "111111111001100111",  "111111111001101010",  "111111111001101101",  "111111111001110000",  "111111111001110011",  "111111111001110110",  "111111111001111001",  "111111111001111100",  "111111111010000000",  "111111111010000011",  "111111111010000110",  "111111111010001001",  "111111111010001100",  "111111111010001111",  "111111111010010010",  "111111111010010101",  "111111111010011000",  "111111111010011011",  "111111111010011110",  "111111111010100010",  "111111111010100101",  "111111111010101000",  "111111111010101011",  "111111111010101110",  "111111111010110001",  "111111111010110100",  "111111111010111000",  "111111111010111011",  "111111111010111110",  "111111111011000001",  "111111111011000100",  "111111111011000111",  "111111111011001011",  "111111111011001110",  "111111111011010001",  "111111111011010100",  "111111111011010111",  "111111111011011010",  "111111111011011110",  "111111111011100001",  "111111111011100100",  "111111111011100111",  "111111111011101010",  "111111111011101110",  "111111111011110001",  "111111111011110100",  "111111111011110111",  "111111111011111011",  "111111111011111110",  "111111111100000001",  "111111111100000100",  "111111111100001000",  "111111111100001011",  "111111111100001110",  "111111111100010001",  "111111111100010101",  "111111111100011000",  "111111111100011011",  "111111111100011110",  "111111111100100010",  "111111111100100101",  "111111111100101000",  "111111111100101100",  "111111111100101111",  "111111111100110010",  "111111111100110101",  "111111111100111001",  "111111111100111100",  "111111111100111111",  "111111111101000011",  "111111111101000110",  "111111111101001001",  "111111111101001101",  "111111111101010000",  "111111111101010011",  "111111111101010111",  "111111111101011010",  "111111111101011101",  "111111111101100001",  "111111111101100100",  "111111111101100111",  "111111111101101011",  "111111111101101110",  "111111111101110001",  "111111111101110101",  "111111111101111000",  "111111111101111011",  "111111111101111111",  "111111111110000010",  "111111111110000101",  "111111111110001001",  "111111111110001100",  "111111111110010000",  "111111111110010011",  "111111111110010110",  "111111111110011010",  "111111111110011101",  "111111111110100000",  "111111111110100100",  "111111111110100111",  "111111111110101011",  "111111111110101110",  "111111111110110001",  "111111111110110101",  "111111111110111000",  "111111111110111100",  "111111111110111111",  "111111111111000010",  "111111111111000110",  "111111111111001001",  "111111111111001101",  "111111111111010000",  "111111111111010011",  "111111111111010111",  "111111111111011010",  "111111111111011110",  "111111111111100001",  "111111111111100101",  "111111111111101000",  "111111111111101011",  "111111111111101111",  "111111111111110010",  "111111111111110110",  "111111111111111001",  "111111111111111101"),("000000000000000000",  "000000000000000011",  "000000000000000111",  "000000000000001010",  "000000000000001110",  "000000000000010001",  "000000000000010101",  "000000000000011000",  "000000000000011100",  "000000000000011111",  "000000000000100010",  "000000000000100110",  "000000000000101001",  "000000000000101101",  "000000000000110000",  "000000000000110100",  "000000000000110111",  "000000000000111011",  "000000000000111110",  "000000000001000001",  "000000000001000101",  "000000000001001000",  "000000000001001100",  "000000000001001111",  "000000000001010011",  "000000000001010110",  "000000000001011010",  "000000000001011101",  "000000000001100001",  "000000000001100100",  "000000000001100111",  "000000000001101011",  "000000000001101110",  "000000000001110010",  "000000000001110101",  "000000000001111001",  "000000000001111100",  "000000000010000000",  "000000000010000011",  "000000000010000111",  "000000000010001010",  "000000000010001110",  "000000000010010001",  "000000000010010100",  "000000000010011000",  "000000000010011011",  "000000000010011111",  "000000000010100010",  "000000000010100110",  "000000000010101001",  "000000000010101101",  "000000000010110000",  "000000000010110100",  "000000000010110111",  "000000000010111011",  "000000000010111110",  "000000000011000001",  "000000000011000101",  "000000000011001000",  "000000000011001100",  "000000000011001111",  "000000000011010011",  "000000000011010110",  "000000000011011010",  "000000000011011101",  "000000000011100001",  "000000000011100100",  "000000000011100111",  "000000000011101011",  "000000000011101110",  "000000000011110010",  "000000000011110101",  "000000000011111001",  "000000000011111100",  "000000000100000000",  "000000000100000011",  "000000000100000110",  "000000000100001010",  "000000000100001101",  "000000000100010001",  "000000000100010100",  "000000000100011000",  "000000000100011011",  "000000000100011110",  "000000000100100010",  "000000000100100101",  "000000000100101001",  "000000000100101100",  "000000000100110000",  "000000000100110011",  "000000000100110110",  "000000000100111010",  "000000000100111101",  "000000000101000001",  "000000000101000100",  "000000000101001000",  "000000000101001011",  "000000000101001110",  "000000000101010010",  "000000000101010101",  "000000000101011001",  "000000000101011100",  "000000000101011111",  "000000000101100011",  "000000000101100110",  "000000000101101010",  "000000000101101101",  "000000000101110000",  "000000000101110100",  "000000000101110111",  "000000000101111010",  "000000000101111110",  "000000000110000001",  "000000000110000101",  "000000000110001000",  "000000000110001011",  "000000000110001111",  "000000000110010010",  "000000000110010101",  "000000000110011001",  "000000000110011100",  "000000000110100000",  "000000000110100011",  "000000000110100110",  "000000000110101010",  "000000000110101101",  "000000000110110000",  "000000000110110100",  "000000000110110111",  "000000000110111010",  "000000000110111110",  "000000000111000001",  "000000000111000100",  "000000000111001000",  "000000000111001011",  "000000000111001110",  "000000000111010010",  "000000000111010101",  "000000000111011000",  "000000000111011011",  "000000000111011111",  "000000000111100010",  "000000000111100101",  "000000000111101001",  "000000000111101100",  "000000000111101111",  "000000000111110010",  "000000000111110110",  "000000000111111001",  "000000000111111100",  "000000001000000000",  "000000001000000011",  "000000001000000110",  "000000001000001001",  "000000001000001101",  "000000001000010000",  "000000001000010011",  "000000001000010110",  "000000001000011010",  "000000001000011101",  "000000001000100000",  "000000001000100011",  "000000001000100110",  "000000001000101010",  "000000001000101101",  "000000001000110000",  "000000001000110011",  "000000001000110110",  "000000001000111010",  "000000001000111101",  "000000001001000000",  "000000001001000011",  "000000001001000110",  "000000001001001010",  "000000001001001101",  "000000001001010000",  "000000001001010011",  "000000001001010110",  "000000001001011001",  "000000001001011101",  "000000001001100000",  "000000001001100011",  "000000001001100110",  "000000001001101001",  "000000001001101100",  "000000001001101111",  "000000001001110010",  "000000001001110110",  "000000001001111001",  "000000001001111100",  "000000001001111111",  "000000001010000010",  "000000001010000101",  "000000001010001000",  "000000001010001011",  "000000001010001110",  "000000001010010001",  "000000001010010100",  "000000001010010111",  "000000001010011011",  "000000001010011110",  "000000001010100001",  "000000001010100100",  "000000001010100111",  "000000001010101010",  "000000001010101101",  "000000001010110000",  "000000001010110011",  "000000001010110110",  "000000001010111001",  "000000001010111100",  "000000001010111111",  "000000001011000010",  "000000001011000101",  "000000001011001000",  "000000001011001011",  "000000001011001110",  "000000001011010001",  "000000001011010011",  "000000001011010110",  "000000001011011001",  "000000001011011100",  "000000001011011111",  "000000001011100010",  "000000001011100101",  "000000001011101000",  "000000001011101011",  "000000001011101110",  "000000001011110001",  "000000001011110100",  "000000001011110110",  "000000001011111001",  "000000001011111100",  "000000001011111111",  "000000001100000010",  "000000001100000101",  "000000001100001000",  "000000001100001010",  "000000001100001101",  "000000001100010000",  "000000001100010011",  "000000001100010110",  "000000001100011000",  "000000001100011011",  "000000001100011110",  "000000001100100001",  "000000001100100100",  "000000001100100110",  "000000001100101001",  "000000001100101100",  "000000001100101111",  "000000001100110001",  "000000001100110100",  "000000001100110111",  "000000001100111010",  "000000001100111100",  "000000001100111111",  "000000001101000010",  "000000001101000100",  "000000001101000111",  "000000001101001010",  "000000001101001100",  "000000001101001111",  "000000001101010010",  "000000001101010100",  "000000001101010111",  "000000001101011010",  "000000001101011100",  "000000001101011111",  "000000001101100010",  "000000001101100100",  "000000001101100111",  "000000001101101001",  "000000001101101100",  "000000001101101111",  "000000001101110001",  "000000001101110100",  "000000001101110110",  "000000001101111001",  "000000001101111011",  "000000001101111110",  "000000001110000000",  "000000001110000011",  "000000001110000110",  "000000001110001000",  "000000001110001011",  "000000001110001101",  "000000001110010000",  "000000001110010010",  "000000001110010100",  "000000001110010111",  "000000001110011001",  "000000001110011100",  "000000001110011110",  "000000001110100001",  "000000001110100011",  "000000001110100110",  "000000001110101000",  "000000001110101010",  "000000001110101101",  "000000001110101111",  "000000001110110001",  "000000001110110100",  "000000001110110110",  "000000001110111001",  "000000001110111011",  "000000001110111101",  "000000001111000000",  "000000001111000010",  "000000001111000100",  "000000001111000111",  "000000001111001001",  "000000001111001011",  "000000001111001101",  "000000001111010000",  "000000001111010010",  "000000001111010100",  "000000001111010110",  "000000001111011001",  "000000001111011011",  "000000001111011101",  "000000001111011111",  "000000001111100001",  "000000001111100100",  "000000001111100110",  "000000001111101000",  "000000001111101010",  "000000001111101100",  "000000001111101111",  "000000001111110001",  "000000001111110011",  "000000001111110101",  "000000001111110111",  "000000001111111001",  "000000001111111011",  "000000001111111101",  "000000001111111111",  "000000010000000001",  "000000010000000100",  "000000010000000110",  "000000010000001000",  "000000010000001010",  "000000010000001100",  "000000010000001110",  "000000010000010000",  "000000010000010010",  "000000010000010100",  "000000010000010110",  "000000010000011000",  "000000010000011010",  "000000010000011100",  "000000010000011110",  "000000010000011111",  "000000010000100001",  "000000010000100011",  "000000010000100101",  "000000010000100111",  "000000010000101001",  "000000010000101011",  "000000010000101101",  "000000010000101111",  "000000010000110000",  "000000010000110010",  "000000010000110100",  "000000010000110110",  "000000010000111000",  "000000010000111010",  "000000010000111011",  "000000010000111101",  "000000010000111111",  "000000010001000001",  "000000010001000010",  "000000010001000100",  "000000010001000110",  "000000010001001000",  "000000010001001001",  "000000010001001011",  "000000010001001101",  "000000010001001110",  "000000010001010000",  "000000010001010010",  "000000010001010011",  "000000010001010101",  "000000010001010111",  "000000010001011000",  "000000010001011010",  "000000010001011100",  "000000010001011101",  "000000010001011111",  "000000010001100000",  "000000010001100010",  "000000010001100100",  "000000010001100101",  "000000010001100111",  "000000010001101000",  "000000010001101010",  "000000010001101011",  "000000010001101101",  "000000010001101110",  "000000010001110000",  "000000010001110001",  "000000010001110011",  "000000010001110100",  "000000010001110101",  "000000010001110111",  "000000010001111000",  "000000010001111010",  "000000010001111011",  "000000010001111100",  "000000010001111110",  "000000010001111111",  "000000010010000001",  "000000010010000010",  "000000010010000011",  "000000010010000101",  "000000010010000110",  "000000010010000111",  "000000010010001000",  "000000010010001010",  "000000010010001011",  "000000010010001100",  "000000010010001110",  "000000010010001111",  "000000010010010000",  "000000010010010001",  "000000010010010010",  "000000010010010100",  "000000010010010101",  "000000010010010110",  "000000010010010111",  "000000010010011000",  "000000010010011001",  "000000010010011011",  "000000010010011100",  "000000010010011101",  "000000010010011110",  "000000010010011111",  "000000010010100000",  "000000010010100001",  "000000010010100010",  "000000010010100011",  "000000010010100100",  "000000010010100101",  "000000010010100110",  "000000010010100111",  "000000010010101000",  "000000010010101001",  "000000010010101010",  "000000010010101011",  "000000010010101100",  "000000010010101101",  "000000010010101110",  "000000010010101111",  "000000010010110000",  "000000010010110001",  "000000010010110010",  "000000010010110011",  "000000010010110011",  "000000010010110100",  "000000010010110101",  "000000010010110110",  "000000010010110111",  "000000010010111000",  "000000010010111000",  "000000010010111001",  "000000010010111010",  "000000010010111011",  "000000010010111011",  "000000010010111100",  "000000010010111101",  "000000010010111110",  "000000010010111110",  "000000010010111111",  "000000010011000000",  "000000010011000000",  "000000010011000001",  "000000010011000010",  "000000010011000010",  "000000010011000011",  "000000010011000100",  "000000010011000100",  "000000010011000101",  "000000010011000101",  "000000010011000110",  "000000010011000110",  "000000010011000111",  "000000010011001000",  "000000010011001000",  "000000010011001001",  "000000010011001001",  "000000010011001010",  "000000010011001010",  "000000010011001010",  "000000010011001011",  "000000010011001011",  "000000010011001100",  "000000010011001100",  "000000010011001101",  "000000010011001101",  "000000010011001101",  "000000010011001110",  "000000010011001110",  "000000010011001111",  "000000010011001111",  "000000010011001111",  "000000010011010000",  "000000010011010000",  "000000010011010000",  "000000010011010000",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010000",  "000000010011010000",  "000000010011010000",  "000000010011001111",  "000000010011001111",  "000000010011001111",  "000000010011001110",  "000000010011001110",  "000000010011001110",  "000000010011001101",  "000000010011001101",  "000000010011001101",  "000000010011001100",  "000000010011001100",  "000000010011001011",  "000000010011001011",  "000000010011001010",  "000000010011001010",  "000000010011001001",  "000000010011001001",  "000000010011001000",  "000000010011001000",  "000000010011000111",  "000000010011000111",  "000000010011000110",  "000000010011000110",  "000000010011000101",  "000000010011000100",  "000000010011000100",  "000000010011000011",  "000000010011000011",  "000000010011000010",  "000000010011000001",  "000000010011000001",  "000000010011000000",  "000000010010111111",  "000000010010111111",  "000000010010111110",  "000000010010111101",  "000000010010111100",  "000000010010111100",  "000000010010111011",  "000000010010111010",  "000000010010111001",  "000000010010111001",  "000000010010111000",  "000000010010110111",  "000000010010110110",  "000000010010110101",  "000000010010110100",  "000000010010110100",  "000000010010110011",  "000000010010110010",  "000000010010110001",  "000000010010110000",  "000000010010101111",  "000000010010101110",  "000000010010101101",  "000000010010101100",  "000000010010101011",  "000000010010101010",  "000000010010101001",  "000000010010101000",  "000000010010100111",  "000000010010100110",  "000000010010100101",  "000000010010100100",  "000000010010100011",  "000000010010100010",  "000000010010100001",  "000000010010100000",  "000000010010011111",  "000000010010011110",  "000000010010011100",  "000000010010011011",  "000000010010011010",  "000000010010011001",  "000000010010011000",  "000000010010010111",  "000000010010010101",  "000000010010010100",  "000000010010010011",  "000000010010010010",  "000000010010010001",  "000000010010001111",  "000000010010001110",  "000000010010001101",  "000000010010001011",  "000000010010001010",  "000000010010001001",  "000000010010000111",  "000000010010000110",  "000000010010000101",  "000000010010000011",  "000000010010000010",  "000000010010000001",  "000000010001111111",  "000000010001111110",  "000000010001111100",  "000000010001111011",  "000000010001111010",  "000000010001111000",  "000000010001110111",  "000000010001110101",  "000000010001110100",  "000000010001110010",  "000000010001110001",  "000000010001101111",  "000000010001101110",  "000000010001101100",  "000000010001101011",  "000000010001101001",  "000000010001100111",  "000000010001100110",  "000000010001100100",  "000000010001100011",  "000000010001100001",  "000000010001011111",  "000000010001011110",  "000000010001011100",  "000000010001011010",  "000000010001011001",  "000000010001010111",  "000000010001010101",  "000000010001010100",  "000000010001010010",  "000000010001010000",  "000000010001001110",  "000000010001001101",  "000000010001001011",  "000000010001001001",  "000000010001000111",  "000000010001000101",  "000000010001000100",  "000000010001000010",  "000000010001000000",  "000000010000111110",  "000000010000111100",  "000000010000111010",  "000000010000111001",  "000000010000110111",  "000000010000110101",  "000000010000110011",  "000000010000110001",  "000000010000101111",  "000000010000101101",  "000000010000101011",  "000000010000101001",  "000000010000100111",  "000000010000100101",  "000000010000100011",  "000000010000100001",  "000000010000011111",  "000000010000011101",  "000000010000011011",  "000000010000011001",  "000000010000010111",  "000000010000010101",  "000000010000010011",  "000000010000010001",  "000000010000001111",  "000000010000001101",  "000000010000001010",  "000000010000001000",  "000000010000000110",  "000000010000000100",  "000000010000000010",  "000000010000000000",  "000000001111111101",  "000000001111111011",  "000000001111111001",  "000000001111110111",  "000000001111110101",  "000000001111110010",  "000000001111110000",  "000000001111101110",  "000000001111101100",  "000000001111101001",  "000000001111100111",  "000000001111100101",  "000000001111100010",  "000000001111100000",  "000000001111011110",  "000000001111011011",  "000000001111011001",  "000000001111010111",  "000000001111010100",  "000000001111010010",  "000000001111001111",  "000000001111001101",  "000000001111001011",  "000000001111001000",  "000000001111000110",  "000000001111000011",  "000000001111000001",  "000000001110111110",  "000000001110111100",  "000000001110111001",  "000000001110110111",  "000000001110110100",  "000000001110110010",  "000000001110101111",  "000000001110101101",  "000000001110101010",  "000000001110101000",  "000000001110100101",  "000000001110100011",  "000000001110100000",  "000000001110011101",  "000000001110011011",  "000000001110011000",  "000000001110010110",  "000000001110010011",  "000000001110010000",  "000000001110001110",  "000000001110001011",  "000000001110001000",  "000000001110000110",  "000000001110000011",  "000000001110000000",  "000000001101111110",  "000000001101111011",  "000000001101111000",  "000000001101110101",  "000000001101110011",  "000000001101110000",  "000000001101101101",  "000000001101101010",  "000000001101101000",  "000000001101100101",  "000000001101100010",  "000000001101011111",  "000000001101011100",  "000000001101011010",  "000000001101010111",  "000000001101010100",  "000000001101010001",  "000000001101001110",  "000000001101001011",  "000000001101001000",  "000000001101000110",  "000000001101000011",  "000000001101000000",  "000000001100111101",  "000000001100111010",  "000000001100110111",  "000000001100110100",  "000000001100110001",  "000000001100101110",  "000000001100101011",  "000000001100101000",  "000000001100100101",  "000000001100100010",  "000000001100011111",  "000000001100011100",  "000000001100011001",  "000000001100010110",  "000000001100010011",  "000000001100010000",  "000000001100001101",  "000000001100001010",  "000000001100000111",  "000000001100000100",  "000000001100000001",  "000000001011111101",  "000000001011111010",  "000000001011110111",  "000000001011110100",  "000000001011110001",  "000000001011101110",  "000000001011101011",  "000000001011100111",  "000000001011100100",  "000000001011100001",  "000000001011011110",  "000000001011011011",  "000000001011011000",  "000000001011010100",  "000000001011010001",  "000000001011001110",  "000000001011001011",  "000000001011000111",  "000000001011000100",  "000000001011000001",  "000000001010111110",  "000000001010111010",  "000000001010110111",  "000000001010110100",  "000000001010110001",  "000000001010101101",  "000000001010101010",  "000000001010100111",  "000000001010100011",  "000000001010100000",  "000000001010011101",  "000000001010011001",  "000000001010010110",  "000000001010010011",  "000000001010001111",  "000000001010001100",  "000000001010001000",  "000000001010000101",  "000000001010000010",  "000000001001111110",  "000000001001111011",  "000000001001110111",  "000000001001110100",  "000000001001110000",  "000000001001101101",  "000000001001101010",  "000000001001100110",  "000000001001100011",  "000000001001011111",  "000000001001011100",  "000000001001011000",  "000000001001010101",  "000000001001010001",  "000000001001001110",  "000000001001001010",  "000000001001000111",  "000000001001000011",  "000000001001000000",  "000000001000111100",  "000000001000111001",  "000000001000110101",  "000000001000110001",  "000000001000101110",  "000000001000101010",  "000000001000100111",  "000000001000100011",  "000000001000011111",  "000000001000011100",  "000000001000011000",  "000000001000010101",  "000000001000010001",  "000000001000001101",  "000000001000001010",  "000000001000000110",  "000000001000000010",  "000000000111111111",  "000000000111111011",  "000000000111110111",  "000000000111110100",  "000000000111110000",  "000000000111101100",  "000000000111101001",  "000000000111100101",  "000000000111100001",  "000000000111011110",  "000000000111011010",  "000000000111010110",  "000000000111010011",  "000000000111001111",  "000000000111001011",  "000000000111000111",  "000000000111000100",  "000000000111000000",  "000000000110111100",  "000000000110111000",  "000000000110110101",  "000000000110110001",  "000000000110101101",  "000000000110101001",  "000000000110100101",  "000000000110100010",  "000000000110011110",  "000000000110011010",  "000000000110010110",  "000000000110010010",  "000000000110001111",  "000000000110001011",  "000000000110000111",  "000000000110000011",  "000000000101111111",  "000000000101111011",  "000000000101110111",  "000000000101110100",  "000000000101110000",  "000000000101101100",  "000000000101101000",  "000000000101100100",  "000000000101100000",  "000000000101011100",  "000000000101011000",  "000000000101010101",  "000000000101010001",  "000000000101001101",  "000000000101001001",  "000000000101000101",  "000000000101000001",  "000000000100111101",  "000000000100111001",  "000000000100110101",  "000000000100110001",  "000000000100101101",  "000000000100101001",  "000000000100100101",  "000000000100100001",  "000000000100011101",  "000000000100011010",  "000000000100010110",  "000000000100010010",  "000000000100001110",  "000000000100001010",  "000000000100000110",  "000000000100000010",  "000000000011111110",  "000000000011111010",  "000000000011110110",  "000000000011110010",  "000000000011101110",  "000000000011101010",  "000000000011100110",  "000000000011100010",  "000000000011011110",  "000000000011011010",  "000000000011010110",  "000000000011010001",  "000000000011001101",  "000000000011001001",  "000000000011000101",  "000000000011000001",  "000000000010111101",  "000000000010111001",  "000000000010110101",  "000000000010110001",  "000000000010101101",  "000000000010101001",  "000000000010100101",  "000000000010100001",  "000000000010011101",  "000000000010011001",  "000000000010010101",  "000000000010010001",  "000000000010001100",  "000000000010001000",  "000000000010000100",  "000000000010000000",  "000000000001111100",  "000000000001111000",  "000000000001110100",  "000000000001110000",  "000000000001101100",  "000000000001101000",  "000000000001100011",  "000000000001011111",  "000000000001011011",  "000000000001010111",  "000000000001010011",  "000000000001001111",  "000000000001001011",  "000000000001000111",  "000000000001000010",  "000000000000111110",  "000000000000111010",  "000000000000110110",  "000000000000110010",  "000000000000101110",  "000000000000101010",  "000000000000100101",  "000000000000100001",  "000000000000011101",  "000000000000011001",  "000000000000010101",  "000000000000010001",  "000000000000001100",  "000000000000001000",  "000000000000000100"),("000000000000000000",  "111111111111111100",  "111111111111111000",  "111111111111110100",  "111111111111101111",  "111111111111101011",  "111111111111100111",  "111111111111100011",  "111111111111011111",  "111111111111011010",  "111111111111010110",  "111111111111010010",  "111111111111001110",  "111111111111001010",  "111111111111000110",  "111111111111000001",  "111111111110111101",  "111111111110111001",  "111111111110110101",  "111111111110110001",  "111111111110101100",  "111111111110101000",  "111111111110100100",  "111111111110100000",  "111111111110011100",  "111111111110011000",  "111111111110010011",  "111111111110001111",  "111111111110001011",  "111111111110000111",  "111111111110000011",  "111111111101111110",  "111111111101111010",  "111111111101110110",  "111111111101110010",  "111111111101101110",  "111111111101101001",  "111111111101100101",  "111111111101100001",  "111111111101011101",  "111111111101011001",  "111111111101010100",  "111111111101010000",  "111111111101001100",  "111111111101001000",  "111111111101000100",  "111111111100111111",  "111111111100111011",  "111111111100110111",  "111111111100110011",  "111111111100101111",  "111111111100101011",  "111111111100100110",  "111111111100100010",  "111111111100011110",  "111111111100011010",  "111111111100010110",  "111111111100010001",  "111111111100001101",  "111111111100001001",  "111111111100000101",  "111111111100000001",  "111111111011111100",  "111111111011111000",  "111111111011110100",  "111111111011110000",  "111111111011101100",  "111111111011101000",  "111111111011100011",  "111111111011011111",  "111111111011011011",  "111111111011010111",  "111111111011010011",  "111111111011001110",  "111111111011001010",  "111111111011000110",  "111111111011000010",  "111111111010111110",  "111111111010111010",  "111111111010110101",  "111111111010110001",  "111111111010101101",  "111111111010101001",  "111111111010100101",  "111111111010100001",  "111111111010011101",  "111111111010011000",  "111111111010010100",  "111111111010010000",  "111111111010001100",  "111111111010001000",  "111111111010000100",  "111111111010000000",  "111111111001111011",  "111111111001110111",  "111111111001110011",  "111111111001101111",  "111111111001101011",  "111111111001100111",  "111111111001100011",  "111111111001011110",  "111111111001011010",  "111111111001010110",  "111111111001010010",  "111111111001001110",  "111111111001001010",  "111111111001000110",  "111111111001000010",  "111111111000111110",  "111111111000111001",  "111111111000110101",  "111111111000110001",  "111111111000101101",  "111111111000101001",  "111111111000100101",  "111111111000100001",  "111111111000011101",  "111111111000011001",  "111111111000010101",  "111111111000010001",  "111111111000001101",  "111111111000001001",  "111111111000000100",  "111111111000000000",  "111111110111111100",  "111111110111111000",  "111111110111110100",  "111111110111110000",  "111111110111101100",  "111111110111101000",  "111111110111100100",  "111111110111100000",  "111111110111011100",  "111111110111011000",  "111111110111010100",  "111111110111010000",  "111111110111001100",  "111111110111001000",  "111111110111000100",  "111111110111000000",  "111111110110111100",  "111111110110111000",  "111111110110110100",  "111111110110110000",  "111111110110101100",  "111111110110101000",  "111111110110100100",  "111111110110100000",  "111111110110011100",  "111111110110011000",  "111111110110010100",  "111111110110010000",  "111111110110001100",  "111111110110001000",  "111111110110000101",  "111111110110000001",  "111111110101111101",  "111111110101111001",  "111111110101110101",  "111111110101110001",  "111111110101101101",  "111111110101101001",  "111111110101100101",  "111111110101100001",  "111111110101011101",  "111111110101011010",  "111111110101010110",  "111111110101010010",  "111111110101001110",  "111111110101001010",  "111111110101000110",  "111111110101000010",  "111111110100111111",  "111111110100111011",  "111111110100110111",  "111111110100110011",  "111111110100101111",  "111111110100101011",  "111111110100101000",  "111111110100100100",  "111111110100100000",  "111111110100011100",  "111111110100011000",  "111111110100010101",  "111111110100010001",  "111111110100001101",  "111111110100001001",  "111111110100000101",  "111111110100000010",  "111111110011111110",  "111111110011111010",  "111111110011110110",  "111111110011110011",  "111111110011101111",  "111111110011101011",  "111111110011101000",  "111111110011100100",  "111111110011100000",  "111111110011011100",  "111111110011011001",  "111111110011010101",  "111111110011010001",  "111111110011001110",  "111111110011001010",  "111111110011000110",  "111111110011000011",  "111111110010111111",  "111111110010111011",  "111111110010111000",  "111111110010110100",  "111111110010110001",  "111111110010101101",  "111111110010101001",  "111111110010100110",  "111111110010100010",  "111111110010011111",  "111111110010011011",  "111111110010010111",  "111111110010010100",  "111111110010010000",  "111111110010001101",  "111111110010001001",  "111111110010000110",  "111111110010000010",  "111111110001111111",  "111111110001111011",  "111111110001111000",  "111111110001110100",  "111111110001110001",  "111111110001101101",  "111111110001101010",  "111111110001100110",  "111111110001100011",  "111111110001011111",  "111111110001011100",  "111111110001011000",  "111111110001010101",  "111111110001010001",  "111111110001001110",  "111111110001001011",  "111111110001000111",  "111111110001000100",  "111111110001000000",  "111111110000111101",  "111111110000111010",  "111111110000110110",  "111111110000110011",  "111111110000110000",  "111111110000101100",  "111111110000101001",  "111111110000100110",  "111111110000100010",  "111111110000011111",  "111111110000011100",  "111111110000011000",  "111111110000010101",  "111111110000010010",  "111111110000001111",  "111111110000001011",  "111111110000001000",  "111111110000000101",  "111111110000000010",  "111111101111111110",  "111111101111111011",  "111111101111111000",  "111111101111110101",  "111111101111110010",  "111111101111101110",  "111111101111101011",  "111111101111101000",  "111111101111100101",  "111111101111100010",  "111111101111011111",  "111111101111011011",  "111111101111011000",  "111111101111010101",  "111111101111010010",  "111111101111001111",  "111111101111001100",  "111111101111001001",  "111111101111000110",  "111111101111000011",  "111111101111000000",  "111111101110111101",  "111111101110111010",  "111111101110110111",  "111111101110110100",  "111111101110110001",  "111111101110101110",  "111111101110101011",  "111111101110101000",  "111111101110100101",  "111111101110100010",  "111111101110011111",  "111111101110011100",  "111111101110011001",  "111111101110010110",  "111111101110010011",  "111111101110010000",  "111111101110001101",  "111111101110001010",  "111111101110001000",  "111111101110000101",  "111111101110000010",  "111111101101111111",  "111111101101111100",  "111111101101111001",  "111111101101110111",  "111111101101110100",  "111111101101110001",  "111111101101101110",  "111111101101101011",  "111111101101101001",  "111111101101100110",  "111111101101100011",  "111111101101100000",  "111111101101011110",  "111111101101011011",  "111111101101011000",  "111111101101010110",  "111111101101010011",  "111111101101010000",  "111111101101001110",  "111111101101001011",  "111111101101001000",  "111111101101000110",  "111111101101000011",  "111111101101000000",  "111111101100111110",  "111111101100111011",  "111111101100111001",  "111111101100110110",  "111111101100110100",  "111111101100110001",  "111111101100101110",  "111111101100101100",  "111111101100101001",  "111111101100100111",  "111111101100100100",  "111111101100100010",  "111111101100100000",  "111111101100011101",  "111111101100011011",  "111111101100011000",  "111111101100010110",  "111111101100010011",  "111111101100010001",  "111111101100001111",  "111111101100001100",  "111111101100001010",  "111111101100000111",  "111111101100000101",  "111111101100000011",  "111111101100000000",  "111111101011111110",  "111111101011111100",  "111111101011111010",  "111111101011110111",  "111111101011110101",  "111111101011110011",  "111111101011110001",  "111111101011101110",  "111111101011101100",  "111111101011101010",  "111111101011101000",  "111111101011100101",  "111111101011100011",  "111111101011100001",  "111111101011011111",  "111111101011011101",  "111111101011011011",  "111111101011011001",  "111111101011010110",  "111111101011010100",  "111111101011010010",  "111111101011010000",  "111111101011001110",  "111111101011001100",  "111111101011001010",  "111111101011001000",  "111111101011000110",  "111111101011000100",  "111111101011000010",  "111111101011000000",  "111111101010111110",  "111111101010111100",  "111111101010111010",  "111111101010111000",  "111111101010110110",  "111111101010110100",  "111111101010110011",  "111111101010110001",  "111111101010101111",  "111111101010101101",  "111111101010101011",  "111111101010101001",  "111111101010101000",  "111111101010100110",  "111111101010100100",  "111111101010100010",  "111111101010100000",  "111111101010011111",  "111111101010011101",  "111111101010011011",  "111111101010011001",  "111111101010011000",  "111111101010010110",  "111111101010010100",  "111111101010010011",  "111111101010010001",  "111111101010001111",  "111111101010001110",  "111111101010001100",  "111111101010001010",  "111111101010001001",  "111111101010000111",  "111111101010000110",  "111111101010000100",  "111111101010000011",  "111111101010000001",  "111111101010000000",  "111111101001111110",  "111111101001111101",  "111111101001111011",  "111111101001111010",  "111111101001111000",  "111111101001110111",  "111111101001110101",  "111111101001110100",  "111111101001110011",  "111111101001110001",  "111111101001110000",  "111111101001101110",  "111111101001101101",  "111111101001101100",  "111111101001101010",  "111111101001101001",  "111111101001101000",  "111111101001100110",  "111111101001100101",  "111111101001100100",  "111111101001100011",  "111111101001100001",  "111111101001100000",  "111111101001011111",  "111111101001011110",  "111111101001011101",  "111111101001011100",  "111111101001011010",  "111111101001011001",  "111111101001011000",  "111111101001010111",  "111111101001010110",  "111111101001010101",  "111111101001010100",  "111111101001010011",  "111111101001010010",  "111111101001010001",  "111111101001010000",  "111111101001001111",  "111111101001001110",  "111111101001001101",  "111111101001001100",  "111111101001001011",  "111111101001001010",  "111111101001001001",  "111111101001001000",  "111111101001000111",  "111111101001000110",  "111111101001000101",  "111111101001000100",  "111111101001000100",  "111111101001000011",  "111111101001000010",  "111111101001000001",  "111111101001000000",  "111111101000111111",  "111111101000111111",  "111111101000111110",  "111111101000111101",  "111111101000111101",  "111111101000111100",  "111111101000111011",  "111111101000111010",  "111111101000111010",  "111111101000111001",  "111111101000111000",  "111111101000111000",  "111111101000110111",  "111111101000110111",  "111111101000110110",  "111111101000110101",  "111111101000110101",  "111111101000110100",  "111111101000110100",  "111111101000110011",  "111111101000110011",  "111111101000110010",  "111111101000110010",  "111111101000110001",  "111111101000110001",  "111111101000110001",  "111111101000110000",  "111111101000110000",  "111111101000101111",  "111111101000101111",  "111111101000101111",  "111111101000101110",  "111111101000101110",  "111111101000101110",  "111111101000101101",  "111111101000101101",  "111111101000101101",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101101",  "111111101000101101",  "111111101000101101",  "111111101000101110",  "111111101000101110",  "111111101000101110",  "111111101000101111",  "111111101000101111",  "111111101000101111",  "111111101000110000",  "111111101000110000",  "111111101000110001",  "111111101000110001",  "111111101000110010",  "111111101000110010",  "111111101000110010",  "111111101000110011",  "111111101000110011",  "111111101000110100",  "111111101000110101",  "111111101000110101",  "111111101000110110",  "111111101000110110",  "111111101000110111",  "111111101000110111",  "111111101000111000",  "111111101000111001",  "111111101000111001",  "111111101000111010",  "111111101000111011",  "111111101000111011",  "111111101000111100",  "111111101000111101",  "111111101000111110",  "111111101000111110",  "111111101000111111",  "111111101001000000",  "111111101001000001",  "111111101001000010",  "111111101001000010",  "111111101001000011",  "111111101001000100",  "111111101001000101",  "111111101001000110",  "111111101001000111",  "111111101001001000",  "111111101001001001",  "111111101001001001",  "111111101001001010",  "111111101001001011",  "111111101001001100",  "111111101001001101",  "111111101001001110",  "111111101001001111",  "111111101001010000",  "111111101001010001",  "111111101001010011",  "111111101001010100",  "111111101001010101",  "111111101001010110",  "111111101001010111",  "111111101001011000",  "111111101001011001",  "111111101001011010",  "111111101001011100",  "111111101001011101",  "111111101001011110",  "111111101001011111",  "111111101001100000",  "111111101001100010",  "111111101001100011",  "111111101001100100",  "111111101001100110",  "111111101001100111",  "111111101001101000",  "111111101001101001",  "111111101001101011",  "111111101001101100",  "111111101001101110",  "111111101001101111",  "111111101001110000",  "111111101001110010",  "111111101001110011",  "111111101001110101",  "111111101001110110",  "111111101001111000",  "111111101001111001",  "111111101001111011",  "111111101001111100",  "111111101001111110",  "111111101001111111",  "111111101010000001",  "111111101010000010",  "111111101010000100",  "111111101010000101",  "111111101010000111",  "111111101010001001",  "111111101010001010",  "111111101010001100",  "111111101010001110",  "111111101010001111",  "111111101010010001",  "111111101010010011",  "111111101010010100",  "111111101010010110",  "111111101010011000",  "111111101010011010",  "111111101010011011",  "111111101010011101",  "111111101010011111",  "111111101010100001",  "111111101010100011",  "111111101010100101",  "111111101010100110",  "111111101010101000",  "111111101010101010",  "111111101010101100",  "111111101010101110",  "111111101010110000",  "111111101010110010",  "111111101010110100",  "111111101010110110",  "111111101010111000",  "111111101010111010",  "111111101010111100",  "111111101010111110",  "111111101011000000",  "111111101011000010",  "111111101011000100",  "111111101011000110",  "111111101011001000",  "111111101011001010",  "111111101011001100",  "111111101011001110",  "111111101011010001",  "111111101011010011",  "111111101011010101",  "111111101011010111",  "111111101011011001",  "111111101011011011",  "111111101011011110",  "111111101011100000",  "111111101011100010",  "111111101011100100",  "111111101011100111",  "111111101011101001",  "111111101011101011",  "111111101011101110",  "111111101011110000",  "111111101011110010",  "111111101011110101",  "111111101011110111",  "111111101011111001",  "111111101011111100",  "111111101011111110",  "111111101100000001",  "111111101100000011",  "111111101100000101",  "111111101100001000",  "111111101100001010",  "111111101100001101",  "111111101100001111",  "111111101100010010",  "111111101100010100",  "111111101100010111",  "111111101100011001",  "111111101100011100",  "111111101100011111",  "111111101100100001",  "111111101100100100",  "111111101100100110",  "111111101100101001",  "111111101100101100",  "111111101100101110",  "111111101100110001",  "111111101100110100",  "111111101100110110",  "111111101100111001",  "111111101100111100",  "111111101100111110",  "111111101101000001",  "111111101101000100",  "111111101101000111",  "111111101101001001",  "111111101101001100",  "111111101101001111",  "111111101101010010",  "111111101101010101",  "111111101101011000",  "111111101101011010",  "111111101101011101",  "111111101101100000",  "111111101101100011",  "111111101101100110",  "111111101101101001",  "111111101101101100",  "111111101101101111",  "111111101101110010",  "111111101101110101",  "111111101101111000",  "111111101101111011",  "111111101101111110",  "111111101110000001",  "111111101110000100",  "111111101110000111",  "111111101110001010",  "111111101110001101",  "111111101110010000",  "111111101110010011",  "111111101110010110",  "111111101110011001",  "111111101110011100",  "111111101110011111",  "111111101110100010",  "111111101110100110",  "111111101110101001",  "111111101110101100",  "111111101110101111",  "111111101110110010",  "111111101110110101",  "111111101110111001",  "111111101110111100",  "111111101110111111",  "111111101111000010",  "111111101111000110",  "111111101111001001",  "111111101111001100",  "111111101111010000",  "111111101111010011",  "111111101111010110",  "111111101111011001",  "111111101111011101",  "111111101111100000",  "111111101111100100",  "111111101111100111",  "111111101111101010",  "111111101111101110",  "111111101111110001",  "111111101111110101",  "111111101111111000",  "111111101111111011",  "111111101111111111",  "111111110000000010",  "111111110000000110",  "111111110000001001",  "111111110000001101",  "111111110000010000",  "111111110000010100",  "111111110000010111",  "111111110000011011",  "111111110000011110",  "111111110000100010",  "111111110000100110",  "111111110000101001",  "111111110000101101",  "111111110000110000",  "111111110000110100",  "111111110000111000",  "111111110000111011",  "111111110000111111",  "111111110001000011",  "111111110001000110",  "111111110001001010",  "111111110001001110",  "111111110001010001",  "111111110001010101",  "111111110001011001",  "111111110001011100",  "111111110001100000",  "111111110001100100",  "111111110001101000",  "111111110001101011",  "111111110001101111",  "111111110001110011",  "111111110001110111",  "111111110001111011",  "111111110001111110",  "111111110010000010",  "111111110010000110",  "111111110010001010",  "111111110010001110",  "111111110010010010",  "111111110010010110",  "111111110010011001",  "111111110010011101",  "111111110010100001",  "111111110010100101",  "111111110010101001",  "111111110010101101",  "111111110010110001",  "111111110010110101",  "111111110010111001",  "111111110010111101",  "111111110011000001",  "111111110011000101",  "111111110011001001",  "111111110011001101",  "111111110011010001",  "111111110011010101",  "111111110011011001",  "111111110011011101",  "111111110011100001",  "111111110011100101",  "111111110011101001",  "111111110011101101",  "111111110011110001",  "111111110011110101",  "111111110011111010",  "111111110011111110",  "111111110100000010",  "111111110100000110",  "111111110100001010",  "111111110100001110",  "111111110100010010",  "111111110100010111",  "111111110100011011",  "111111110100011111",  "111111110100100011",  "111111110100100111",  "111111110100101100",  "111111110100110000",  "111111110100110100",  "111111110100111000",  "111111110100111101",  "111111110101000001",  "111111110101000101",  "111111110101001001",  "111111110101001110",  "111111110101010010",  "111111110101010110",  "111111110101011010",  "111111110101011111",  "111111110101100011",  "111111110101100111",  "111111110101101100",  "111111110101110000",  "111111110101110100",  "111111110101111001",  "111111110101111101",  "111111110110000010",  "111111110110000110",  "111111110110001010",  "111111110110001111",  "111111110110010011",  "111111110110011000",  "111111110110011100",  "111111110110100000",  "111111110110100101",  "111111110110101001",  "111111110110101110",  "111111110110110010",  "111111110110110111",  "111111110110111011",  "111111110111000000",  "111111110111000100",  "111111110111001001",  "111111110111001101",  "111111110111010010",  "111111110111010110",  "111111110111011011",  "111111110111011111",  "111111110111100100",  "111111110111101000",  "111111110111101101",  "111111110111110001",  "111111110111110110",  "111111110111111010",  "111111110111111111",  "111111111000000100",  "111111111000001000",  "111111111000001101",  "111111111000010001",  "111111111000010110",  "111111111000011011",  "111111111000011111",  "111111111000100100",  "111111111000101000",  "111111111000101101",  "111111111000110010",  "111111111000110110",  "111111111000111011",  "111111111001000000",  "111111111001000100",  "111111111001001001",  "111111111001001110",  "111111111001010010",  "111111111001010111",  "111111111001011100",  "111111111001100000",  "111111111001100101",  "111111111001101010",  "111111111001101111",  "111111111001110011",  "111111111001111000",  "111111111001111101",  "111111111010000001",  "111111111010000110",  "111111111010001011",  "111111111010010000",  "111111111010010100",  "111111111010011001",  "111111111010011110",  "111111111010100011",  "111111111010101000",  "111111111010101100",  "111111111010110001",  "111111111010110110",  "111111111010111011",  "111111111011000000",  "111111111011000100",  "111111111011001001",  "111111111011001110",  "111111111011010011",  "111111111011011000",  "111111111011011100",  "111111111011100001",  "111111111011100110",  "111111111011101011",  "111111111011110000",  "111111111011110101",  "111111111011111010",  "111111111011111110",  "111111111100000011",  "111111111100001000",  "111111111100001101",  "111111111100010010",  "111111111100010111",  "111111111100011100",  "111111111100100001",  "111111111100100101",  "111111111100101010",  "111111111100101111",  "111111111100110100",  "111111111100111001",  "111111111100111110",  "111111111101000011",  "111111111101001000",  "111111111101001101",  "111111111101010010",  "111111111101010111",  "111111111101011100",  "111111111101100000",  "111111111101100101",  "111111111101101010",  "111111111101101111",  "111111111101110100",  "111111111101111001",  "111111111101111110",  "111111111110000011",  "111111111110001000",  "111111111110001101",  "111111111110010010",  "111111111110010111",  "111111111110011100",  "111111111110100001",  "111111111110100110",  "111111111110101011",  "111111111110110000",  "111111111110110101",  "111111111110111010",  "111111111110111111",  "111111111111000100",  "111111111111001001",  "111111111111001110",  "111111111111010011",  "111111111111011000",  "111111111111011101",  "111111111111100010",  "111111111111100111",  "111111111111101100",  "111111111111110001",  "111111111111110110",  "111111111111111011"),("000000000000000000",  "000000000000000101",  "000000000000001010",  "000000000000001111",  "000000000000010100",  "000000000000011001",  "000000000000011110",  "000000000000100011",  "000000000000101000",  "000000000000101101",  "000000000000110010",  "000000000000110111",  "000000000000111100",  "000000000001000001",  "000000000001000110",  "000000000001001100",  "000000000001010001",  "000000000001010110",  "000000000001011011",  "000000000001100000",  "000000000001100101",  "000000000001101010",  "000000000001101111",  "000000000001110100",  "000000000001111001",  "000000000001111110",  "000000000010000011",  "000000000010001000",  "000000000010001101",  "000000000010010010",  "000000000010010111",  "000000000010011100",  "000000000010100001",  "000000000010100110",  "000000000010101011",  "000000000010110001",  "000000000010110110",  "000000000010111011",  "000000000011000000",  "000000000011000101",  "000000000011001010",  "000000000011001111",  "000000000011010100",  "000000000011011001",  "000000000011011110",  "000000000011100011",  "000000000011101000",  "000000000011101101",  "000000000011110010",  "000000000011110111",  "000000000011111100",  "000000000100000001",  "000000000100000110",  "000000000100001100",  "000000000100010001",  "000000000100010110",  "000000000100011011",  "000000000100100000",  "000000000100100101",  "000000000100101010",  "000000000100101111",  "000000000100110100",  "000000000100111001",  "000000000100111110",  "000000000101000011",  "000000000101001000",  "000000000101001101",  "000000000101010010",  "000000000101010111",  "000000000101011100",  "000000000101100001",  "000000000101100110",  "000000000101101011",  "000000000101110000",  "000000000101110101",  "000000000101111010",  "000000000101111111",  "000000000110000100",  "000000000110001001",  "000000000110001111",  "000000000110010100",  "000000000110011001",  "000000000110011110",  "000000000110100011",  "000000000110101000",  "000000000110101101",  "000000000110110010",  "000000000110110111",  "000000000110111100",  "000000000111000001",  "000000000111000110",  "000000000111001011",  "000000000111010000",  "000000000111010101",  "000000000111011010",  "000000000111011111",  "000000000111100011",  "000000000111101000",  "000000000111101101",  "000000000111110010",  "000000000111110111",  "000000000111111100",  "000000001000000001",  "000000001000000110",  "000000001000001011",  "000000001000010000",  "000000001000010101",  "000000001000011010",  "000000001000011111",  "000000001000100100",  "000000001000101001",  "000000001000101110",  "000000001000110011",  "000000001000111000",  "000000001000111101",  "000000001001000001",  "000000001001000110",  "000000001001001011",  "000000001001010000",  "000000001001010101",  "000000001001011010",  "000000001001011111",  "000000001001100100",  "000000001001101001",  "000000001001101110",  "000000001001110010",  "000000001001110111",  "000000001001111100",  "000000001010000001",  "000000001010000110",  "000000001010001011",  "000000001010010000",  "000000001010010100",  "000000001010011001",  "000000001010011110",  "000000001010100011",  "000000001010101000",  "000000001010101101",  "000000001010110001",  "000000001010110110",  "000000001010111011",  "000000001011000000",  "000000001011000101",  "000000001011001010",  "000000001011001110",  "000000001011010011",  "000000001011011000",  "000000001011011101",  "000000001011100001",  "000000001011100110",  "000000001011101011",  "000000001011110000",  "000000001011110100",  "000000001011111001",  "000000001011111110",  "000000001100000011",  "000000001100000111",  "000000001100001100",  "000000001100010001",  "000000001100010110",  "000000001100011010",  "000000001100011111",  "000000001100100100",  "000000001100101000",  "000000001100101101",  "000000001100110010",  "000000001100110110",  "000000001100111011",  "000000001101000000",  "000000001101000100",  "000000001101001001",  "000000001101001110",  "000000001101010010",  "000000001101010111",  "000000001101011011",  "000000001101100000",  "000000001101100101",  "000000001101101001",  "000000001101101110",  "000000001101110010",  "000000001101110111",  "000000001101111100",  "000000001110000000",  "000000001110000101",  "000000001110001001",  "000000001110001110",  "000000001110010010",  "000000001110010111",  "000000001110011011",  "000000001110100000",  "000000001110100100",  "000000001110101001",  "000000001110101101",  "000000001110110010",  "000000001110110110",  "000000001110111011",  "000000001110111111",  "000000001111000100",  "000000001111001000",  "000000001111001101",  "000000001111010001",  "000000001111010110",  "000000001111011010",  "000000001111011110",  "000000001111100011",  "000000001111100111",  "000000001111101100",  "000000001111110000",  "000000001111110100",  "000000001111111001",  "000000001111111101",  "000000010000000001",  "000000010000000110",  "000000010000001010",  "000000010000001110",  "000000010000010011",  "000000010000010111",  "000000010000011011",  "000000010000100000",  "000000010000100100",  "000000010000101000",  "000000010000101101",  "000000010000110001",  "000000010000110101",  "000000010000111001",  "000000010000111110",  "000000010001000010",  "000000010001000110",  "000000010001001010",  "000000010001001110",  "000000010001010011",  "000000010001010111",  "000000010001011011",  "000000010001011111",  "000000010001100011",  "000000010001100111",  "000000010001101011",  "000000010001110000",  "000000010001110100",  "000000010001111000",  "000000010001111100",  "000000010010000000",  "000000010010000100",  "000000010010001000",  "000000010010001100",  "000000010010010000",  "000000010010010100",  "000000010010011000",  "000000010010011100",  "000000010010100000",  "000000010010100100",  "000000010010101000",  "000000010010101100",  "000000010010110000",  "000000010010110100",  "000000010010111000",  "000000010010111100",  "000000010011000000",  "000000010011000100",  "000000010011001000",  "000000010011001100",  "000000010011010000",  "000000010011010100",  "000000010011010111",  "000000010011011011",  "000000010011011111",  "000000010011100011",  "000000010011100111",  "000000010011101011",  "000000010011101110",  "000000010011110010",  "000000010011110110",  "000000010011111010",  "000000010011111110",  "000000010100000001",  "000000010100000101",  "000000010100001001",  "000000010100001101",  "000000010100010000",  "000000010100010100",  "000000010100011000",  "000000010100011011",  "000000010100011111",  "000000010100100011",  "000000010100100110",  "000000010100101010",  "000000010100101110",  "000000010100110001",  "000000010100110101",  "000000010100111000",  "000000010100111100",  "000000010101000000",  "000000010101000011",  "000000010101000111",  "000000010101001010",  "000000010101001110",  "000000010101010001",  "000000010101010101",  "000000010101011000",  "000000010101011100",  "000000010101011111",  "000000010101100011",  "000000010101100110",  "000000010101101001",  "000000010101101101",  "000000010101110000",  "000000010101110100",  "000000010101110111",  "000000010101111010",  "000000010101111110",  "000000010110000001",  "000000010110000100",  "000000010110001000",  "000000010110001011",  "000000010110001110",  "000000010110010010",  "000000010110010101",  "000000010110011000",  "000000010110011011",  "000000010110011111",  "000000010110100010",  "000000010110100101",  "000000010110101000",  "000000010110101011",  "000000010110101111",  "000000010110110010",  "000000010110110101",  "000000010110111000",  "000000010110111011",  "000000010110111110",  "000000010111000001",  "000000010111000100",  "000000010111001000",  "000000010111001011",  "000000010111001110",  "000000010111010001",  "000000010111010100",  "000000010111010111",  "000000010111011010",  "000000010111011101",  "000000010111100000",  "000000010111100011",  "000000010111100110",  "000000010111101000",  "000000010111101011",  "000000010111101110",  "000000010111110001",  "000000010111110100",  "000000010111110111",  "000000010111111010",  "000000010111111101",  "000000010111111111",  "000000011000000010",  "000000011000000101",  "000000011000001000",  "000000011000001011",  "000000011000001101",  "000000011000010000",  "000000011000010011",  "000000011000010101",  "000000011000011000",  "000000011000011011",  "000000011000011101",  "000000011000100000",  "000000011000100011",  "000000011000100101",  "000000011000101000",  "000000011000101011",  "000000011000101101",  "000000011000110000",  "000000011000110010",  "000000011000110101",  "000000011000110111",  "000000011000111010",  "000000011000111100",  "000000011000111111",  "000000011001000001",  "000000011001000100",  "000000011001000110",  "000000011001001001",  "000000011001001011",  "000000011001001110",  "000000011001010000",  "000000011001010010",  "000000011001010101",  "000000011001010111",  "000000011001011001",  "000000011001011100",  "000000011001011110",  "000000011001100000",  "000000011001100010",  "000000011001100101",  "000000011001100111",  "000000011001101001",  "000000011001101011",  "000000011001101110",  "000000011001110000",  "000000011001110010",  "000000011001110100",  "000000011001110110",  "000000011001111000",  "000000011001111010",  "000000011001111101",  "000000011001111111",  "000000011010000001",  "000000011010000011",  "000000011010000101",  "000000011010000111",  "000000011010001001",  "000000011010001011",  "000000011010001101",  "000000011010001111",  "000000011010010001",  "000000011010010011",  "000000011010010101",  "000000011010010110",  "000000011010011000",  "000000011010011010",  "000000011010011100",  "000000011010011110",  "000000011010100000",  "000000011010100001",  "000000011010100011",  "000000011010100101",  "000000011010100111",  "000000011010101001",  "000000011010101010",  "000000011010101100",  "000000011010101110",  "000000011010101111",  "000000011010110001",  "000000011010110011",  "000000011010110100",  "000000011010110110",  "000000011010111000",  "000000011010111001",  "000000011010111011",  "000000011010111100",  "000000011010111110",  "000000011010111111",  "000000011011000001",  "000000011011000010",  "000000011011000100",  "000000011011000101",  "000000011011000111",  "000000011011001000",  "000000011011001010",  "000000011011001011",  "000000011011001100",  "000000011011001110",  "000000011011001111",  "000000011011010000",  "000000011011010010",  "000000011011010011",  "000000011011010100",  "000000011011010110",  "000000011011010111",  "000000011011011000",  "000000011011011001",  "000000011011011010",  "000000011011011100",  "000000011011011101",  "000000011011011110",  "000000011011011111",  "000000011011100000",  "000000011011100001",  "000000011011100010",  "000000011011100100",  "000000011011100101",  "000000011011100110",  "000000011011100111",  "000000011011101000",  "000000011011101001",  "000000011011101010",  "000000011011101011",  "000000011011101100",  "000000011011101100",  "000000011011101101",  "000000011011101110",  "000000011011101111",  "000000011011110000",  "000000011011110001",  "000000011011110010",  "000000011011110011",  "000000011011110011",  "000000011011110100",  "000000011011110101",  "000000011011110110",  "000000011011110110",  "000000011011110111",  "000000011011111000",  "000000011011111000",  "000000011011111001",  "000000011011111010",  "000000011011111010",  "000000011011111011",  "000000011011111100",  "000000011011111100",  "000000011011111101",  "000000011011111101",  "000000011011111110",  "000000011011111110",  "000000011011111111",  "000000011011111111",  "000000011100000000",  "000000011100000000",  "000000011100000001",  "000000011100000001",  "000000011100000001",  "000000011100000010",  "000000011100000010",  "000000011100000011",  "000000011100000011",  "000000011100000011",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000011",  "000000011100000011",  "000000011100000011",  "000000011100000010",  "000000011100000010",  "000000011100000001",  "000000011100000001",  "000000011100000001",  "000000011100000000",  "000000011100000000",  "000000011011111111",  "000000011011111111",  "000000011011111110",  "000000011011111110",  "000000011011111101",  "000000011011111101",  "000000011011111100",  "000000011011111100",  "000000011011111011",  "000000011011111010",  "000000011011111010",  "000000011011111001",  "000000011011111000",  "000000011011111000",  "000000011011110111",  "000000011011110110",  "000000011011110101",  "000000011011110101",  "000000011011110100",  "000000011011110011",  "000000011011110010",  "000000011011110001",  "000000011011110001",  "000000011011110000",  "000000011011101111",  "000000011011101110",  "000000011011101101",  "000000011011101100",  "000000011011101011",  "000000011011101010",  "000000011011101001",  "000000011011101000",  "000000011011100111",  "000000011011100110",  "000000011011100101",  "000000011011100100",  "000000011011100011",  "000000011011100010",  "000000011011100001",  "000000011011100000",  "000000011011011111",  "000000011011011101",  "000000011011011100",  "000000011011011011",  "000000011011011010",  "000000011011011001",  "000000011011010111",  "000000011011010110",  "000000011011010101",  "000000011011010011",  "000000011011010010",  "000000011011010001",  "000000011011001111",  "000000011011001110",  "000000011011001101",  "000000011011001011",  "000000011011001010",  "000000011011001000",  "000000011011000111",  "000000011011000101",  "000000011011000100",  "000000011011000010",  "000000011011000001",  "000000011010111111",  "000000011010111110",  "000000011010111100",  "000000011010111011",  "000000011010111001",  "000000011010110111",  "000000011010110110",  "000000011010110100",  "000000011010110010",  "000000011010110001",  "000000011010101111",  "000000011010101101",  "000000011010101100",  "000000011010101010",  "000000011010101000",  "000000011010100110",  "000000011010100100",  "000000011010100011",  "000000011010100001",  "000000011010011111",  "000000011010011101",  "000000011010011011",  "000000011010011001",  "000000011010010111",  "000000011010010101",  "000000011010010011",  "000000011010010001",  "000000011010001111",  "000000011010001101",  "000000011010001011",  "000000011010001001",  "000000011010000111",  "000000011010000101",  "000000011010000011",  "000000011010000001",  "000000011001111111",  "000000011001111101",  "000000011001111010",  "000000011001111000",  "000000011001110110",  "000000011001110100",  "000000011001110010",  "000000011001101111",  "000000011001101101",  "000000011001101011",  "000000011001101001",  "000000011001100110",  "000000011001100100",  "000000011001100010",  "000000011001011111",  "000000011001011101",  "000000011001011011",  "000000011001011000",  "000000011001010110",  "000000011001010011",  "000000011001010001",  "000000011001001110",  "000000011001001100",  "000000011001001001",  "000000011001000111",  "000000011001000100",  "000000011001000010",  "000000011000111111",  "000000011000111101",  "000000011000111010",  "000000011000110111",  "000000011000110101",  "000000011000110010",  "000000011000101111",  "000000011000101101",  "000000011000101010",  "000000011000100111",  "000000011000100101",  "000000011000100010",  "000000011000011111",  "000000011000011100",  "000000011000011010",  "000000011000010111",  "000000011000010100",  "000000011000010001",  "000000011000001110",  "000000011000001011",  "000000011000001001",  "000000011000000110",  "000000011000000011",  "000000011000000000",  "000000010111111101",  "000000010111111010",  "000000010111110111",  "000000010111110100",  "000000010111110001",  "000000010111101110",  "000000010111101011",  "000000010111101000",  "000000010111100101",  "000000010111100010",  "000000010111011111",  "000000010111011011",  "000000010111011000",  "000000010111010101",  "000000010111010010",  "000000010111001111",  "000000010111001100",  "000000010111001000",  "000000010111000101",  "000000010111000010",  "000000010110111111",  "000000010110111011",  "000000010110111000",  "000000010110110101",  "000000010110110010",  "000000010110101110",  "000000010110101011",  "000000010110101000",  "000000010110100100",  "000000010110100001",  "000000010110011101",  "000000010110011010",  "000000010110010111",  "000000010110010011",  "000000010110010000",  "000000010110001100",  "000000010110001001",  "000000010110000101",  "000000010110000010",  "000000010101111110",  "000000010101111011",  "000000010101110111",  "000000010101110011",  "000000010101110000",  "000000010101101100",  "000000010101101001",  "000000010101100101",  "000000010101100001",  "000000010101011110",  "000000010101011010",  "000000010101010110",  "000000010101010011",  "000000010101001111",  "000000010101001011",  "000000010101000111",  "000000010101000100",  "000000010101000000",  "000000010100111100",  "000000010100111000",  "000000010100110100",  "000000010100110001",  "000000010100101101",  "000000010100101001",  "000000010100100101",  "000000010100100001",  "000000010100011101",  "000000010100011001",  "000000010100010101",  "000000010100010001",  "000000010100001110",  "000000010100001010",  "000000010100000110",  "000000010100000010",  "000000010011111110",  "000000010011111010",  "000000010011110101",  "000000010011110001",  "000000010011101101",  "000000010011101001",  "000000010011100101",  "000000010011100001",  "000000010011011101",  "000000010011011001",  "000000010011010101",  "000000010011010001",  "000000010011001100",  "000000010011001000",  "000000010011000100",  "000000010011000000",  "000000010010111100",  "000000010010110111",  "000000010010110011",  "000000010010101111",  "000000010010101011",  "000000010010100110",  "000000010010100010",  "000000010010011110",  "000000010010011001",  "000000010010010101",  "000000010010010001",  "000000010010001100",  "000000010010001000",  "000000010010000100",  "000000010001111111",  "000000010001111011",  "000000010001110110",  "000000010001110010",  "000000010001101101",  "000000010001101001",  "000000010001100100",  "000000010001100000",  "000000010001011011",  "000000010001010111",  "000000010001010010",  "000000010001001110",  "000000010001001001",  "000000010001000101",  "000000010001000000",  "000000010000111100",  "000000010000110111",  "000000010000110010",  "000000010000101110",  "000000010000101001",  "000000010000100101",  "000000010000100000",  "000000010000011011",  "000000010000010111",  "000000010000010010",  "000000010000001101",  "000000010000001000",  "000000010000000100",  "000000001111111111",  "000000001111111010",  "000000001111110101",  "000000001111110001",  "000000001111101100",  "000000001111100111",  "000000001111100010",  "000000001111011110",  "000000001111011001",  "000000001111010100",  "000000001111001111",  "000000001111001010",  "000000001111000101",  "000000001111000000",  "000000001110111100",  "000000001110110111",  "000000001110110010",  "000000001110101101",  "000000001110101000",  "000000001110100011",  "000000001110011110",  "000000001110011001",  "000000001110010100",  "000000001110001111",  "000000001110001010",  "000000001110000101",  "000000001110000000",  "000000001101111011",  "000000001101110110",  "000000001101110001",  "000000001101101100",  "000000001101100111",  "000000001101100010",  "000000001101011101",  "000000001101011000",  "000000001101010010",  "000000001101001101",  "000000001101001000",  "000000001101000011",  "000000001100111110",  "000000001100111001",  "000000001100110100",  "000000001100101110",  "000000001100101001",  "000000001100100100",  "000000001100011111",  "000000001100011010",  "000000001100010100",  "000000001100001111",  "000000001100001010",  "000000001100000101",  "000000001011111111",  "000000001011111010",  "000000001011110101",  "000000001011110000",  "000000001011101010",  "000000001011100101",  "000000001011100000",  "000000001011011010",  "000000001011010101",  "000000001011010000",  "000000001011001010",  "000000001011000101",  "000000001011000000",  "000000001010111010",  "000000001010110101",  "000000001010101111",  "000000001010101010",  "000000001010100101",  "000000001010011111",  "000000001010011010",  "000000001010010100",  "000000001010001111",  "000000001010001001",  "000000001010000100",  "000000001001111111",  "000000001001111001",  "000000001001110100",  "000000001001101110",  "000000001001101001",  "000000001001100011",  "000000001001011110",  "000000001001011000",  "000000001001010011",  "000000001001001101",  "000000001001000111",  "000000001001000010",  "000000001000111100",  "000000001000110111",  "000000001000110001",  "000000001000101100",  "000000001000100110",  "000000001000100000",  "000000001000011011",  "000000001000010101",  "000000001000010000",  "000000001000001010",  "000000001000000100",  "000000000111111111",  "000000000111111001",  "000000000111110011",  "000000000111101110",  "000000000111101000",  "000000000111100010",  "000000000111011101",  "000000000111010111",  "000000000111010001",  "000000000111001100",  "000000000111000110",  "000000000111000000",  "000000000110111011",  "000000000110110101",  "000000000110101111",  "000000000110101001",  "000000000110100100",  "000000000110011110",  "000000000110011000",  "000000000110010010",  "000000000110001101",  "000000000110000111",  "000000000110000001",  "000000000101111011",  "000000000101110110",  "000000000101110000",  "000000000101101010",  "000000000101100100",  "000000000101011110",  "000000000101011001",  "000000000101010011",  "000000000101001101",  "000000000101000111",  "000000000101000001",  "000000000100111011",  "000000000100110110",  "000000000100110000",  "000000000100101010",  "000000000100100100",  "000000000100011110",  "000000000100011000",  "000000000100010010",  "000000000100001100",  "000000000100000111",  "000000000100000001",  "000000000011111011",  "000000000011110101",  "000000000011101111",  "000000000011101001",  "000000000011100011",  "000000000011011101",  "000000000011010111",  "000000000011010001",  "000000000011001100",  "000000000011000110",  "000000000011000000",  "000000000010111010",  "000000000010110100",  "000000000010101110",  "000000000010101000",  "000000000010100010",  "000000000010011100",  "000000000010010110",  "000000000010010000",  "000000000010001010",  "000000000010000100",  "000000000001111110",  "000000000001111000",  "000000000001110010",  "000000000001101100",  "000000000001100110",  "000000000001100000",  "000000000001011010",  "000000000001010100",  "000000000001001110",  "000000000001001000",  "000000000001000010",  "000000000000111100",  "000000000000110110",  "000000000000110000",  "000000000000101010",  "000000000000100100",  "000000000000011110",  "000000000000011000",  "000000000000010010",  "000000000000001100",  "000000000000000110"),("000000000000000000",  "111111111111111010",  "111111111111110100",  "111111111111101110",  "111111111111101000",  "111111111111100010",  "111111111111011100",  "111111111111010110",  "111111111111010000",  "111111111111001010",  "111111111111000100",  "111111111110111110",  "111111111110110111",  "111111111110110001",  "111111111110101011",  "111111111110100101",  "111111111110011111",  "111111111110011001",  "111111111110010011",  "111111111110001101",  "111111111110000111",  "111111111110000001",  "111111111101111011",  "111111111101110101",  "111111111101101111",  "111111111101101001",  "111111111101100011",  "111111111101011101",  "111111111101010110",  "111111111101010000",  "111111111101001010",  "111111111101000100",  "111111111100111110",  "111111111100111000",  "111111111100110010",  "111111111100101100",  "111111111100100110",  "111111111100100000",  "111111111100011010",  "111111111100010100",  "111111111100001110",  "111111111100000111",  "111111111100000001",  "111111111011111011",  "111111111011110101",  "111111111011101111",  "111111111011101001",  "111111111011100011",  "111111111011011101",  "111111111011010111",  "111111111011010001",  "111111111011001011",  "111111111011000101",  "111111111010111111",  "111111111010111001",  "111111111010110010",  "111111111010101100",  "111111111010100110",  "111111111010100000",  "111111111010011010",  "111111111010010100",  "111111111010001110",  "111111111010001000",  "111111111010000010",  "111111111001111100",  "111111111001110110",  "111111111001110000",  "111111111001101010",  "111111111001100100",  "111111111001011110",  "111111111001011000",  "111111111001010010",  "111111111001001100",  "111111111001000110",  "111111111000111111",  "111111111000111001",  "111111111000110011",  "111111111000101101",  "111111111000100111",  "111111111000100001",  "111111111000011011",  "111111111000010101",  "111111111000001111",  "111111111000001001",  "111111111000000011",  "111111110111111101",  "111111110111110111",  "111111110111110001",  "111111110111101011",  "111111110111100101",  "111111110111011111",  "111111110111011001",  "111111110111010011",  "111111110111001101",  "111111110111000111",  "111111110111000001",  "111111110110111011",  "111111110110110101",  "111111110110101111",  "111111110110101001",  "111111110110100011",  "111111110110011101",  "111111110110011000",  "111111110110010010",  "111111110110001100",  "111111110110000110",  "111111110110000000",  "111111110101111010",  "111111110101110100",  "111111110101101110",  "111111110101101000",  "111111110101100010",  "111111110101011100",  "111111110101010110",  "111111110101010000",  "111111110101001010",  "111111110101000101",  "111111110100111111",  "111111110100111001",  "111111110100110011",  "111111110100101101",  "111111110100100111",  "111111110100100001",  "111111110100011011",  "111111110100010110",  "111111110100010000",  "111111110100001010",  "111111110100000100",  "111111110011111110",  "111111110011111000",  "111111110011110010",  "111111110011101101",  "111111110011100111",  "111111110011100001",  "111111110011011011",  "111111110011010101",  "111111110011010000",  "111111110011001010",  "111111110011000100",  "111111110010111110",  "111111110010111000",  "111111110010110011",  "111111110010101101",  "111111110010100111",  "111111110010100001",  "111111110010011100",  "111111110010010110",  "111111110010010000",  "111111110010001010",  "111111110010000101",  "111111110001111111",  "111111110001111001",  "111111110001110100",  "111111110001101110",  "111111110001101000",  "111111110001100011",  "111111110001011101",  "111111110001010111",  "111111110001010010",  "111111110001001100",  "111111110001000110",  "111111110001000001",  "111111110000111011",  "111111110000110101",  "111111110000110000",  "111111110000101010",  "111111110000100101",  "111111110000011111",  "111111110000011001",  "111111110000010100",  "111111110000001110",  "111111110000001001",  "111111110000000011",  "111111101111111101",  "111111101111111000",  "111111101111110010",  "111111101111101101",  "111111101111100111",  "111111101111100010",  "111111101111011100",  "111111101111010111",  "111111101111010001",  "111111101111001100",  "111111101111000110",  "111111101111000001",  "111111101110111011",  "111111101110110110",  "111111101110110001",  "111111101110101011",  "111111101110100110",  "111111101110100000",  "111111101110011011",  "111111101110010110",  "111111101110010000",  "111111101110001011",  "111111101110000101",  "111111101110000000",  "111111101101111011",  "111111101101110101",  "111111101101110000",  "111111101101101011",  "111111101101100101",  "111111101101100000",  "111111101101011011",  "111111101101010101",  "111111101101010000",  "111111101101001011",  "111111101101000110",  "111111101101000000",  "111111101100111011",  "111111101100110110",  "111111101100110001",  "111111101100101100",  "111111101100100110",  "111111101100100001",  "111111101100011100",  "111111101100010111",  "111111101100010010",  "111111101100001100",  "111111101100000111",  "111111101100000010",  "111111101011111101",  "111111101011111000",  "111111101011110011",  "111111101011101110",  "111111101011101001",  "111111101011100100",  "111111101011011111",  "111111101011011010",  "111111101011010101",  "111111101011010000",  "111111101011001010",  "111111101011000101",  "111111101011000000",  "111111101010111100",  "111111101010110111",  "111111101010110010",  "111111101010101101",  "111111101010101000",  "111111101010100011",  "111111101010011110",  "111111101010011001",  "111111101010010100",  "111111101010001111",  "111111101010001010",  "111111101010000101",  "111111101010000001",  "111111101001111100",  "111111101001110111",  "111111101001110010",  "111111101001101101",  "111111101001101001",  "111111101001100100",  "111111101001011111",  "111111101001011010",  "111111101001010110",  "111111101001010001",  "111111101001001100",  "111111101001000111",  "111111101001000011",  "111111101000111110",  "111111101000111001",  "111111101000110101",  "111111101000110000",  "111111101000101011",  "111111101000100111",  "111111101000100010",  "111111101000011110",  "111111101000011001",  "111111101000010100",  "111111101000010000",  "111111101000001011",  "111111101000000111",  "111111101000000010",  "111111100111111110",  "111111100111111001",  "111111100111110101",  "111111100111110000",  "111111100111101100",  "111111100111100111",  "111111100111100011",  "111111100111011111",  "111111100111011010",  "111111100111010110",  "111111100111010001",  "111111100111001101",  "111111100111001001",  "111111100111000100",  "111111100111000000",  "111111100110111100",  "111111100110111000",  "111111100110110011",  "111111100110101111",  "111111100110101011",  "111111100110100110",  "111111100110100010",  "111111100110011110",  "111111100110011010",  "111111100110010110",  "111111100110010010",  "111111100110001101",  "111111100110001001",  "111111100110000101",  "111111100110000001",  "111111100101111101",  "111111100101111001",  "111111100101110101",  "111111100101110001",  "111111100101101101",  "111111100101101001",  "111111100101100101",  "111111100101100001",  "111111100101011101",  "111111100101011001",  "111111100101010101",  "111111100101010001",  "111111100101001101",  "111111100101001001",  "111111100101000101",  "111111100101000001",  "111111100100111101",  "111111100100111001",  "111111100100110110",  "111111100100110010",  "111111100100101110",  "111111100100101010",  "111111100100100110",  "111111100100100011",  "111111100100011111",  "111111100100011011",  "111111100100011000",  "111111100100010100",  "111111100100010000",  "111111100100001101",  "111111100100001001",  "111111100100000101",  "111111100100000010",  "111111100011111110",  "111111100011111010",  "111111100011110111",  "111111100011110011",  "111111100011110000",  "111111100011101100",  "111111100011101001",  "111111100011100101",  "111111100011100010",  "111111100011011110",  "111111100011011011",  "111111100011010111",  "111111100011010100",  "111111100011010001",  "111111100011001101",  "111111100011001010",  "111111100011000111",  "111111100011000011",  "111111100011000000",  "111111100010111101",  "111111100010111001",  "111111100010110110",  "111111100010110011",  "111111100010110000",  "111111100010101100",  "111111100010101001",  "111111100010100110",  "111111100010100011",  "111111100010100000",  "111111100010011101",  "111111100010011001",  "111111100010010110",  "111111100010010011",  "111111100010010000",  "111111100010001101",  "111111100010001010",  "111111100010000111",  "111111100010000100",  "111111100010000001",  "111111100001111110",  "111111100001111011",  "111111100001111000",  "111111100001110101",  "111111100001110010",  "111111100001110000",  "111111100001101101",  "111111100001101010",  "111111100001100111",  "111111100001100100",  "111111100001100001",  "111111100001011111",  "111111100001011100",  "111111100001011001",  "111111100001010111",  "111111100001010100",  "111111100001010001",  "111111100001001110",  "111111100001001100",  "111111100001001001",  "111111100001000111",  "111111100001000100",  "111111100001000001",  "111111100000111111",  "111111100000111100",  "111111100000111010",  "111111100000110111",  "111111100000110101",  "111111100000110010",  "111111100000110000",  "111111100000101101",  "111111100000101011",  "111111100000101001",  "111111100000100110",  "111111100000100100",  "111111100000100010",  "111111100000011111",  "111111100000011101",  "111111100000011011",  "111111100000011000",  "111111100000010110",  "111111100000010100",  "111111100000010010",  "111111100000001111",  "111111100000001101",  "111111100000001011",  "111111100000001001",  "111111100000000111",  "111111100000000101",  "111111100000000011",  "111111100000000001",  "111111011111111110",  "111111011111111100",  "111111011111111010",  "111111011111111000",  "111111011111110110",  "111111011111110101",  "111111011111110011",  "111111011111110001",  "111111011111101111",  "111111011111101101",  "111111011111101011",  "111111011111101001",  "111111011111100111",  "111111011111100110",  "111111011111100100",  "111111011111100010",  "111111011111100000",  "111111011111011111",  "111111011111011101",  "111111011111011011",  "111111011111011001",  "111111011111011000",  "111111011111010110",  "111111011111010101",  "111111011111010011",  "111111011111010001",  "111111011111010000",  "111111011111001110",  "111111011111001101",  "111111011111001011",  "111111011111001010",  "111111011111001000",  "111111011111000111",  "111111011111000101",  "111111011111000100",  "111111011111000011",  "111111011111000001",  "111111011111000000",  "111111011110111111",  "111111011110111101",  "111111011110111100",  "111111011110111011",  "111111011110111010",  "111111011110111000",  "111111011110110111",  "111111011110110110",  "111111011110110101",  "111111011110110100",  "111111011110110010",  "111111011110110001",  "111111011110110000",  "111111011110101111",  "111111011110101110",  "111111011110101101",  "111111011110101100",  "111111011110101011",  "111111011110101010",  "111111011110101001",  "111111011110101000",  "111111011110100111",  "111111011110100110",  "111111011110100110",  "111111011110100101",  "111111011110100100",  "111111011110100011",  "111111011110100010",  "111111011110100010",  "111111011110100001",  "111111011110100000",  "111111011110011111",  "111111011110011111",  "111111011110011110",  "111111011110011101",  "111111011110011101",  "111111011110011100",  "111111011110011011",  "111111011110011011",  "111111011110011010",  "111111011110011010",  "111111011110011001",  "111111011110011001",  "111111011110011000",  "111111011110011000",  "111111011110010111",  "111111011110010111",  "111111011110010111",  "111111011110010110",  "111111011110010110",  "111111011110010110",  "111111011110010101",  "111111011110010101",  "111111011110010101",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010101",  "111111011110010101",  "111111011110010101",  "111111011110010101",  "111111011110010110",  "111111011110010110",  "111111011110010110",  "111111011110010111",  "111111011110010111",  "111111011110011000",  "111111011110011000",  "111111011110011001",  "111111011110011001",  "111111011110011010",  "111111011110011010",  "111111011110011011",  "111111011110011011",  "111111011110011100",  "111111011110011100",  "111111011110011101",  "111111011110011110",  "111111011110011110",  "111111011110011111",  "111111011110100000",  "111111011110100001",  "111111011110100001",  "111111011110100010",  "111111011110100011",  "111111011110100100",  "111111011110100100",  "111111011110100101",  "111111011110100110",  "111111011110100111",  "111111011110101000",  "111111011110101001",  "111111011110101010",  "111111011110101011",  "111111011110101100",  "111111011110101101",  "111111011110101110",  "111111011110101111",  "111111011110110000",  "111111011110110001",  "111111011110110010",  "111111011110110011",  "111111011110110101",  "111111011110110110",  "111111011110110111",  "111111011110111000",  "111111011110111001",  "111111011110111011",  "111111011110111100",  "111111011110111101",  "111111011110111111",  "111111011111000000",  "111111011111000001",  "111111011111000011",  "111111011111000100",  "111111011111000110",  "111111011111000111",  "111111011111001000",  "111111011111001010",  "111111011111001011",  "111111011111001101",  "111111011111001111",  "111111011111010000",  "111111011111010010",  "111111011111010011",  "111111011111010101",  "111111011111010111",  "111111011111011000",  "111111011111011010",  "111111011111011100",  "111111011111011101",  "111111011111011111",  "111111011111100001",  "111111011111100011",  "111111011111100101",  "111111011111100110",  "111111011111101000",  "111111011111101010",  "111111011111101100",  "111111011111101110",  "111111011111110000",  "111111011111110010",  "111111011111110100",  "111111011111110110",  "111111011111111000",  "111111011111111010",  "111111011111111100",  "111111011111111110",  "111111100000000000",  "111111100000000010",  "111111100000000100",  "111111100000000110",  "111111100000001001",  "111111100000001011",  "111111100000001101",  "111111100000001111",  "111111100000010010",  "111111100000010100",  "111111100000010110",  "111111100000011000",  "111111100000011011",  "111111100000011101",  "111111100000100000",  "111111100000100010",  "111111100000100100",  "111111100000100111",  "111111100000101001",  "111111100000101100",  "111111100000101110",  "111111100000110001",  "111111100000110011",  "111111100000110110",  "111111100000111000",  "111111100000111011",  "111111100000111110",  "111111100001000000",  "111111100001000011",  "111111100001000110",  "111111100001001000",  "111111100001001011",  "111111100001001110",  "111111100001010000",  "111111100001010011",  "111111100001010110",  "111111100001011001",  "111111100001011100",  "111111100001011110",  "111111100001100001",  "111111100001100100",  "111111100001100111",  "111111100001101010",  "111111100001101101",  "111111100001110000",  "111111100001110011",  "111111100001110110",  "111111100001111001",  "111111100001111100",  "111111100001111111",  "111111100010000010",  "111111100010000101",  "111111100010001000",  "111111100010001100",  "111111100010001111",  "111111100010010010",  "111111100010010101",  "111111100010011000",  "111111100010011100",  "111111100010011111",  "111111100010100010",  "111111100010100101",  "111111100010101001",  "111111100010101100",  "111111100010101111",  "111111100010110011",  "111111100010110110",  "111111100010111001",  "111111100010111101",  "111111100011000000",  "111111100011000100",  "111111100011000111",  "111111100011001011",  "111111100011001110",  "111111100011010010",  "111111100011010101",  "111111100011011001",  "111111100011011101",  "111111100011100000",  "111111100011100100",  "111111100011100111",  "111111100011101011",  "111111100011101111",  "111111100011110011",  "111111100011110110",  "111111100011111010",  "111111100011111110",  "111111100100000001",  "111111100100000101",  "111111100100001001",  "111111100100001101",  "111111100100010001",  "111111100100010101",  "111111100100011001",  "111111100100011100",  "111111100100100000",  "111111100100100100",  "111111100100101000",  "111111100100101100",  "111111100100110000",  "111111100100110100",  "111111100100111000",  "111111100100111100",  "111111100101000000",  "111111100101000100",  "111111100101001001",  "111111100101001101",  "111111100101010001",  "111111100101010101",  "111111100101011001",  "111111100101011101",  "111111100101100010",  "111111100101100110",  "111111100101101010",  "111111100101101110",  "111111100101110011",  "111111100101110111",  "111111100101111011",  "111111100101111111",  "111111100110000100",  "111111100110001000",  "111111100110001101",  "111111100110010001",  "111111100110010101",  "111111100110011010",  "111111100110011110",  "111111100110100011",  "111111100110100111",  "111111100110101100",  "111111100110110000",  "111111100110110101",  "111111100110111001",  "111111100110111110",  "111111100111000010",  "111111100111000111",  "111111100111001100",  "111111100111010000",  "111111100111010101",  "111111100111011010",  "111111100111011110",  "111111100111100011",  "111111100111101000",  "111111100111101100",  "111111100111110001",  "111111100111110110",  "111111100111111011",  "111111100111111111",  "111111101000000100",  "111111101000001001",  "111111101000001110",  "111111101000010011",  "111111101000011000",  "111111101000011101",  "111111101000100001",  "111111101000100110",  "111111101000101011",  "111111101000110000",  "111111101000110101",  "111111101000111010",  "111111101000111111",  "111111101001000100",  "111111101001001001",  "111111101001001110",  "111111101001010011",  "111111101001011000",  "111111101001011110",  "111111101001100011",  "111111101001101000",  "111111101001101101",  "111111101001110010",  "111111101001110111",  "111111101001111100",  "111111101010000010",  "111111101010000111",  "111111101010001100",  "111111101010010001",  "111111101010010111",  "111111101010011100",  "111111101010100001",  "111111101010100111",  "111111101010101100",  "111111101010110001",  "111111101010110111",  "111111101010111100",  "111111101011000001",  "111111101011000111",  "111111101011001100",  "111111101011010010",  "111111101011010111",  "111111101011011100",  "111111101011100010",  "111111101011100111",  "111111101011101101",  "111111101011110010",  "111111101011111000",  "111111101011111101",  "111111101100000011",  "111111101100001001",  "111111101100001110",  "111111101100010100",  "111111101100011001",  "111111101100011111",  "111111101100100101",  "111111101100101010",  "111111101100110000",  "111111101100110110",  "111111101100111011",  "111111101101000001",  "111111101101000111",  "111111101101001100",  "111111101101010010",  "111111101101011000",  "111111101101011110",  "111111101101100100",  "111111101101101001",  "111111101101101111",  "111111101101110101",  "111111101101111011",  "111111101110000001",  "111111101110000111",  "111111101110001100",  "111111101110010010",  "111111101110011000",  "111111101110011110",  "111111101110100100",  "111111101110101010",  "111111101110110000",  "111111101110110110",  "111111101110111100",  "111111101111000010",  "111111101111001000",  "111111101111001110",  "111111101111010100",  "111111101111011010",  "111111101111100000",  "111111101111100110",  "111111101111101100",  "111111101111110010",  "111111101111111000",  "111111101111111110",  "111111110000000101",  "111111110000001011",  "111111110000010001",  "111111110000010111",  "111111110000011101",  "111111110000100011",  "111111110000101010",  "111111110000110000",  "111111110000110110",  "111111110000111100",  "111111110001000010",  "111111110001001001",  "111111110001001111",  "111111110001010101",  "111111110001011100",  "111111110001100010",  "111111110001101000",  "111111110001101110",  "111111110001110101",  "111111110001111011",  "111111110010000001",  "111111110010001000",  "111111110010001110",  "111111110010010101",  "111111110010011011",  "111111110010100001",  "111111110010101000",  "111111110010101110",  "111111110010110101",  "111111110010111011",  "111111110011000010",  "111111110011001000",  "111111110011001110",  "111111110011010101",  "111111110011011011",  "111111110011100010",  "111111110011101000",  "111111110011101111",  "111111110011110110",  "111111110011111100",  "111111110100000011",  "111111110100001001",  "111111110100010000",  "111111110100010110",  "111111110100011101",  "111111110100100100",  "111111110100101010",  "111111110100110001",  "111111110100110111",  "111111110100111110",  "111111110101000101",  "111111110101001011",  "111111110101010010",  "111111110101011001",  "111111110101011111",  "111111110101100110",  "111111110101101101",  "111111110101110011",  "111111110101111010",  "111111110110000001",  "111111110110001000",  "111111110110001110",  "111111110110010101",  "111111110110011100",  "111111110110100011",  "111111110110101001",  "111111110110110000",  "111111110110110111",  "111111110110111110",  "111111110111000101",  "111111110111001011",  "111111110111010010",  "111111110111011001",  "111111110111100000",  "111111110111100111",  "111111110111101110",  "111111110111110100",  "111111110111111011",  "111111111000000010",  "111111111000001001",  "111111111000010000",  "111111111000010111",  "111111111000011110",  "111111111000100101",  "111111111000101100",  "111111111000110010",  "111111111000111001",  "111111111001000000",  "111111111001000111",  "111111111001001110",  "111111111001010101",  "111111111001011100",  "111111111001100011",  "111111111001101010",  "111111111001110001",  "111111111001111000",  "111111111001111111",  "111111111010000110",  "111111111010001101",  "111111111010010100",  "111111111010011011",  "111111111010100010",  "111111111010101001",  "111111111010110000",  "111111111010110111",  "111111111010111110",  "111111111011000101",  "111111111011001100",  "111111111011010011",  "111111111011011010",  "111111111011100010",  "111111111011101001",  "111111111011110000",  "111111111011110111",  "111111111011111110",  "111111111100000101",  "111111111100001100",  "111111111100010011",  "111111111100011010",  "111111111100100001",  "111111111100101001",  "111111111100110000",  "111111111100110111",  "111111111100111110",  "111111111101000101",  "111111111101001100",  "111111111101010011",  "111111111101011011",  "111111111101100010",  "111111111101101001",  "111111111101110000",  "111111111101110111",  "111111111101111110",  "111111111110000110",  "111111111110001101",  "111111111110010100",  "111111111110011011",  "111111111110100010",  "111111111110101001",  "111111111110110001",  "111111111110111000",  "111111111110111111",  "111111111111000110",  "111111111111001101",  "111111111111010101",  "111111111111011100",  "111111111111100011",  "111111111111101010",  "111111111111110010",  "111111111111111001"),("000000000000000000",  "000000000000000111",  "000000000000001110",  "000000000000010110",  "000000000000011101",  "000000000000100100",  "000000000000101011",  "000000000000110011",  "000000000000111010",  "000000000001000001",  "000000000001001000",  "000000000001010000",  "000000000001010111",  "000000000001011110",  "000000000001100101",  "000000000001101101",  "000000000001110100",  "000000000001111011",  "000000000010000010",  "000000000010001010",  "000000000010010001",  "000000000010011000",  "000000000010100000",  "000000000010100111",  "000000000010101110",  "000000000010110101",  "000000000010111101",  "000000000011000100",  "000000000011001011",  "000000000011010010",  "000000000011011010",  "000000000011100001",  "000000000011101000",  "000000000011110000",  "000000000011110111",  "000000000011111110",  "000000000100000101",  "000000000100001101",  "000000000100010100",  "000000000100011011",  "000000000100100011",  "000000000100101010",  "000000000100110001",  "000000000100111000",  "000000000101000000",  "000000000101000111",  "000000000101001110",  "000000000101010101",  "000000000101011101",  "000000000101100100",  "000000000101101011",  "000000000101110011",  "000000000101111010",  "000000000110000001",  "000000000110001000",  "000000000110010000",  "000000000110010111",  "000000000110011110",  "000000000110100101",  "000000000110101101",  "000000000110110100",  "000000000110111011",  "000000000111000010",  "000000000111001010",  "000000000111010001",  "000000000111011000",  "000000000111100000",  "000000000111100111",  "000000000111101110",  "000000000111110101",  "000000000111111100",  "000000001000000100",  "000000001000001011",  "000000001000010010",  "000000001000011001",  "000000001000100001",  "000000001000101000",  "000000001000101111",  "000000001000110110",  "000000001000111110",  "000000001001000101",  "000000001001001100",  "000000001001010011",  "000000001001011010",  "000000001001100010",  "000000001001101001",  "000000001001110000",  "000000001001110111",  "000000001001111110",  "000000001010000110",  "000000001010001101",  "000000001010010100",  "000000001010011011",  "000000001010100010",  "000000001010101001",  "000000001010110001",  "000000001010111000",  "000000001010111111",  "000000001011000110",  "000000001011001101",  "000000001011010100",  "000000001011011100",  "000000001011100011",  "000000001011101010",  "000000001011110001",  "000000001011111000",  "000000001011111111",  "000000001100000110",  "000000001100001101",  "000000001100010101",  "000000001100011100",  "000000001100100011",  "000000001100101010",  "000000001100110001",  "000000001100111000",  "000000001100111111",  "000000001101000110",  "000000001101001101",  "000000001101010100",  "000000001101011011",  "000000001101100010",  "000000001101101001",  "000000001101110000",  "000000001101110111",  "000000001101111110",  "000000001110000101",  "000000001110001100",  "000000001110010011",  "000000001110011010",  "000000001110100001",  "000000001110101000",  "000000001110101111",  "000000001110110110",  "000000001110111101",  "000000001111000100",  "000000001111001011",  "000000001111010010",  "000000001111011001",  "000000001111100000",  "000000001111100111",  "000000001111101110",  "000000001111110101",  "000000001111111100",  "000000010000000011",  "000000010000001010",  "000000010000010000",  "000000010000010111",  "000000010000011110",  "000000010000100101",  "000000010000101100",  "000000010000110011",  "000000010000111010",  "000000010001000000",  "000000010001000111",  "000000010001001110",  "000000010001010101",  "000000010001011100",  "000000010001100010",  "000000010001101001",  "000000010001110000",  "000000010001110111",  "000000010001111101",  "000000010010000100",  "000000010010001011",  "000000010010010010",  "000000010010011000",  "000000010010011111",  "000000010010100110",  "000000010010101101",  "000000010010110011",  "000000010010111010",  "000000010011000001",  "000000010011000111",  "000000010011001110",  "000000010011010101",  "000000010011011011",  "000000010011100010",  "000000010011101000",  "000000010011101111",  "000000010011110110",  "000000010011111100",  "000000010100000011",  "000000010100001001",  "000000010100010000",  "000000010100010110",  "000000010100011101",  "000000010100100011",  "000000010100101010",  "000000010100110000",  "000000010100110111",  "000000010100111101",  "000000010101000100",  "000000010101001010",  "000000010101010001",  "000000010101010111",  "000000010101011110",  "000000010101100100",  "000000010101101011",  "000000010101110001",  "000000010101110111",  "000000010101111110",  "000000010110000100",  "000000010110001010",  "000000010110010001",  "000000010110010111",  "000000010110011101",  "000000010110100100",  "000000010110101010",  "000000010110110000",  "000000010110110111",  "000000010110111101",  "000000010111000011",  "000000010111001001",  "000000010111010000",  "000000010111010110",  "000000010111011100",  "000000010111100010",  "000000010111101000",  "000000010111101111",  "000000010111110101",  "000000010111111011",  "000000011000000001",  "000000011000000111",  "000000011000001101",  "000000011000010011",  "000000011000011001",  "000000011000011111",  "000000011000100101",  "000000011000101100",  "000000011000110010",  "000000011000111000",  "000000011000111110",  "000000011001000100",  "000000011001001010",  "000000011001010000",  "000000011001010101",  "000000011001011011",  "000000011001100001",  "000000011001100111",  "000000011001101101",  "000000011001110011",  "000000011001111001",  "000000011001111111",  "000000011010000101",  "000000011010001010",  "000000011010010000",  "000000011010010110",  "000000011010011100",  "000000011010100010",  "000000011010100111",  "000000011010101101",  "000000011010110011",  "000000011010111001",  "000000011010111110",  "000000011011000100",  "000000011011001010",  "000000011011001111",  "000000011011010101",  "000000011011011011",  "000000011011100000",  "000000011011100110",  "000000011011101011",  "000000011011110001",  "000000011011110111",  "000000011011111100",  "000000011100000010",  "000000011100000111",  "000000011100001101",  "000000011100010010",  "000000011100011000",  "000000011100011101",  "000000011100100011",  "000000011100101000",  "000000011100101101",  "000000011100110011",  "000000011100111000",  "000000011100111101",  "000000011101000011",  "000000011101001000",  "000000011101001101",  "000000011101010011",  "000000011101011000",  "000000011101011101",  "000000011101100011",  "000000011101101000",  "000000011101101101",  "000000011101110010",  "000000011101110111",  "000000011101111101",  "000000011110000010",  "000000011110000111",  "000000011110001100",  "000000011110010001",  "000000011110010110",  "000000011110011011",  "000000011110100000",  "000000011110100101",  "000000011110101010",  "000000011110101111",  "000000011110110100",  "000000011110111001",  "000000011110111110",  "000000011111000011",  "000000011111001000",  "000000011111001101",  "000000011111010010",  "000000011111010111",  "000000011111011100",  "000000011111100001",  "000000011111100101",  "000000011111101010",  "000000011111101111",  "000000011111110100",  "000000011111111000",  "000000011111111101",  "000000100000000010",  "000000100000000111",  "000000100000001011",  "000000100000010000",  "000000100000010101",  "000000100000011001",  "000000100000011110",  "000000100000100010",  "000000100000100111",  "000000100000101011",  "000000100000110000",  "000000100000110101",  "000000100000111001",  "000000100000111110",  "000000100001000010",  "000000100001000110",  "000000100001001011",  "000000100001001111",  "000000100001010100",  "000000100001011000",  "000000100001011100",  "000000100001100001",  "000000100001100101",  "000000100001101001",  "000000100001101110",  "000000100001110010",  "000000100001110110",  "000000100001111010",  "000000100001111110",  "000000100010000011",  "000000100010000111",  "000000100010001011",  "000000100010001111",  "000000100010010011",  "000000100010010111",  "000000100010011011",  "000000100010011111",  "000000100010100011",  "000000100010100111",  "000000100010101011",  "000000100010101111",  "000000100010110011",  "000000100010110111",  "000000100010111011",  "000000100010111111",  "000000100011000011",  "000000100011000111",  "000000100011001011",  "000000100011001110",  "000000100011010010",  "000000100011010110",  "000000100011011010",  "000000100011011101",  "000000100011100001",  "000000100011100101",  "000000100011101000",  "000000100011101100",  "000000100011110000",  "000000100011110011",  "000000100011110111",  "000000100011111010",  "000000100011111110",  "000000100100000010",  "000000100100000101",  "000000100100001001",  "000000100100001100",  "000000100100001111",  "000000100100010011",  "000000100100010110",  "000000100100011010",  "000000100100011101",  "000000100100100000",  "000000100100100100",  "000000100100100111",  "000000100100101010",  "000000100100101110",  "000000100100110001",  "000000100100110100",  "000000100100110111",  "000000100100111010",  "000000100100111101",  "000000100101000001",  "000000100101000100",  "000000100101000111",  "000000100101001010",  "000000100101001101",  "000000100101010000",  "000000100101010011",  "000000100101010110",  "000000100101011001",  "000000100101011100",  "000000100101011111",  "000000100101100010",  "000000100101100100",  "000000100101100111",  "000000100101101010",  "000000100101101101",  "000000100101110000",  "000000100101110010",  "000000100101110101",  "000000100101111000",  "000000100101111011",  "000000100101111101",  "000000100110000000",  "000000100110000011",  "000000100110000101",  "000000100110001000",  "000000100110001010",  "000000100110001101",  "000000100110001111",  "000000100110010010",  "000000100110010100",  "000000100110010111",  "000000100110011001",  "000000100110011100",  "000000100110011110",  "000000100110100000",  "000000100110100011",  "000000100110100101",  "000000100110100111",  "000000100110101010",  "000000100110101100",  "000000100110101110",  "000000100110110000",  "000000100110110011",  "000000100110110101",  "000000100110110111",  "000000100110111001",  "000000100110111011",  "000000100110111101",  "000000100110111111",  "000000100111000001",  "000000100111000011",  "000000100111000101",  "000000100111000111",  "000000100111001001",  "000000100111001011",  "000000100111001101",  "000000100111001111",  "000000100111010001",  "000000100111010010",  "000000100111010100",  "000000100111010110",  "000000100111011000",  "000000100111011001",  "000000100111011011",  "000000100111011101",  "000000100111011110",  "000000100111100000",  "000000100111100010",  "000000100111100011",  "000000100111100101",  "000000100111100110",  "000000100111101000",  "000000100111101001",  "000000100111101011",  "000000100111101100",  "000000100111101110",  "000000100111101111",  "000000100111110000",  "000000100111110010",  "000000100111110011",  "000000100111110100",  "000000100111110110",  "000000100111110111",  "000000100111111000",  "000000100111111001",  "000000100111111011",  "000000100111111100",  "000000100111111101",  "000000100111111110",  "000000100111111111",  "000000101000000000",  "000000101000000001",  "000000101000000010",  "000000101000000011",  "000000101000000100",  "000000101000000101",  "000000101000000110",  "000000101000000111",  "000000101000001000",  "000000101000001001",  "000000101000001001",  "000000101000001010",  "000000101000001011",  "000000101000001100",  "000000101000001101",  "000000101000001101",  "000000101000001110",  "000000101000001111",  "000000101000001111",  "000000101000010000",  "000000101000010000",  "000000101000010001",  "000000101000010010",  "000000101000010010",  "000000101000010011",  "000000101000010011",  "000000101000010011",  "000000101000010100",  "000000101000010100",  "000000101000010101",  "000000101000010101",  "000000101000010101",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010101",  "000000101000010101",  "000000101000010101",  "000000101000010100",  "000000101000010100",  "000000101000010100",  "000000101000010011",  "000000101000010011",  "000000101000010010",  "000000101000010010",  "000000101000010001",  "000000101000010001",  "000000101000010000",  "000000101000001111",  "000000101000001111",  "000000101000001110",  "000000101000001101",  "000000101000001101",  "000000101000001100",  "000000101000001011",  "000000101000001010",  "000000101000001010",  "000000101000001001",  "000000101000001000",  "000000101000000111",  "000000101000000110",  "000000101000000101",  "000000101000000100",  "000000101000000011",  "000000101000000010",  "000000101000000001",  "000000101000000000",  "000000100111111111",  "000000100111111110",  "000000100111111101",  "000000100111111100",  "000000100111111011",  "000000100111111001",  "000000100111111000",  "000000100111110111",  "000000100111110110",  "000000100111110100",  "000000100111110011",  "000000100111110010",  "000000100111110000",  "000000100111101111",  "000000100111101110",  "000000100111101100",  "000000100111101011",  "000000100111101001",  "000000100111101000",  "000000100111100110",  "000000100111100101",  "000000100111100011",  "000000100111100001",  "000000100111100000",  "000000100111011110",  "000000100111011100",  "000000100111011011",  "000000100111011001",  "000000100111010111",  "000000100111010101",  "000000100111010100",  "000000100111010010",  "000000100111010000",  "000000100111001110",  "000000100111001100",  "000000100111001010",  "000000100111001000",  "000000100111000110",  "000000100111000100",  "000000100111000010",  "000000100111000000",  "000000100110111110",  "000000100110111100",  "000000100110111010",  "000000100110111000",  "000000100110110110",  "000000100110110011",  "000000100110110001",  "000000100110101111",  "000000100110101101",  "000000100110101010",  "000000100110101000",  "000000100110100110",  "000000100110100011",  "000000100110100001",  "000000100110011110",  "000000100110011100",  "000000100110011010",  "000000100110010111",  "000000100110010101",  "000000100110010010",  "000000100110001111",  "000000100110001101",  "000000100110001010",  "000000100110001000",  "000000100110000101",  "000000100110000010",  "000000100110000000",  "000000100101111101",  "000000100101111010",  "000000100101110111",  "000000100101110101",  "000000100101110010",  "000000100101101111",  "000000100101101100",  "000000100101101001",  "000000100101100110",  "000000100101100011",  "000000100101100000",  "000000100101011101",  "000000100101011010",  "000000100101010111",  "000000100101010100",  "000000100101010001",  "000000100101001110",  "000000100101001011",  "000000100101001000",  "000000100101000100",  "000000100101000001",  "000000100100111110",  "000000100100111011",  "000000100100111000",  "000000100100110100",  "000000100100110001",  "000000100100101110",  "000000100100101010",  "000000100100100111",  "000000100100100011",  "000000100100100000",  "000000100100011101",  "000000100100011001",  "000000100100010110",  "000000100100010010",  "000000100100001110",  "000000100100001011",  "000000100100000111",  "000000100100000100",  "000000100100000000",  "000000100011111100",  "000000100011111001",  "000000100011110101",  "000000100011110001",  "000000100011101101",  "000000100011101010",  "000000100011100110",  "000000100011100010",  "000000100011011110",  "000000100011011010",  "000000100011010110",  "000000100011010010",  "000000100011001111",  "000000100011001011",  "000000100011000111",  "000000100011000011",  "000000100010111111",  "000000100010111010",  "000000100010110110",  "000000100010110010",  "000000100010101110",  "000000100010101010",  "000000100010100110",  "000000100010100010",  "000000100010011101",  "000000100010011001",  "000000100010010101",  "000000100010010001",  "000000100010001100",  "000000100010001000",  "000000100010000100",  "000000100001111111",  "000000100001111011",  "000000100001110111",  "000000100001110010",  "000000100001101110",  "000000100001101001",  "000000100001100101",  "000000100001100000",  "000000100001011100",  "000000100001010111",  "000000100001010010",  "000000100001001110",  "000000100001001001",  "000000100001000101",  "000000100001000000",  "000000100000111011",  "000000100000110110",  "000000100000110010",  "000000100000101101",  "000000100000101000",  "000000100000100011",  "000000100000011111",  "000000100000011010",  "000000100000010101",  "000000100000010000",  "000000100000001011",  "000000100000000110",  "000000100000000001",  "000000011111111100",  "000000011111110111",  "000000011111110010",  "000000011111101101",  "000000011111101000",  "000000011111100011",  "000000011111011110",  "000000011111011001",  "000000011111010100",  "000000011111001111",  "000000011111001001",  "000000011111000100",  "000000011110111111",  "000000011110111010",  "000000011110110100",  "000000011110101111",  "000000011110101010",  "000000011110100100",  "000000011110011111",  "000000011110011010",  "000000011110010100",  "000000011110001111",  "000000011110001010",  "000000011110000100",  "000000011101111111",  "000000011101111001",  "000000011101110100",  "000000011101101110",  "000000011101101001",  "000000011101100011",  "000000011101011101",  "000000011101011000",  "000000011101010010",  "000000011101001101",  "000000011101000111",  "000000011101000001",  "000000011100111011",  "000000011100110110",  "000000011100110000",  "000000011100101010",  "000000011100100100",  "000000011100011111",  "000000011100011001",  "000000011100010011",  "000000011100001101",  "000000011100000111",  "000000011100000001",  "000000011011111011",  "000000011011110110",  "000000011011110000",  "000000011011101010",  "000000011011100100",  "000000011011011110",  "000000011011011000",  "000000011011010010",  "000000011011001011",  "000000011011000101",  "000000011010111111",  "000000011010111001",  "000000011010110011",  "000000011010101101",  "000000011010100111",  "000000011010100000",  "000000011010011010",  "000000011010010100",  "000000011010001110",  "000000011010001000",  "000000011010000001",  "000000011001111011",  "000000011001110101",  "000000011001101110",  "000000011001101000",  "000000011001100010",  "000000011001011011",  "000000011001010101",  "000000011001001110",  "000000011001001000",  "000000011001000001",  "000000011000111011",  "000000011000110100",  "000000011000101110",  "000000011000100111",  "000000011000100001",  "000000011000011010",  "000000011000010100",  "000000011000001101",  "000000011000000110",  "000000011000000000",  "000000010111111001",  "000000010111110010",  "000000010111101100",  "000000010111100101",  "000000010111011110",  "000000010111011000",  "000000010111010001",  "000000010111001010",  "000000010111000011",  "000000010110111101",  "000000010110110110",  "000000010110101111",  "000000010110101000",  "000000010110100001",  "000000010110011010",  "000000010110010011",  "000000010110001100",  "000000010110000110",  "000000010101111111",  "000000010101111000",  "000000010101110001",  "000000010101101010",  "000000010101100011",  "000000010101011100",  "000000010101010101",  "000000010101001110",  "000000010101000111",  "000000010100111111",  "000000010100111000",  "000000010100110001",  "000000010100101010",  "000000010100100011",  "000000010100011100",  "000000010100010101",  "000000010100001101",  "000000010100000110",  "000000010011111111",  "000000010011111000",  "000000010011110001",  "000000010011101001",  "000000010011100010",  "000000010011011011",  "000000010011010011",  "000000010011001100",  "000000010011000101",  "000000010010111101",  "000000010010110110",  "000000010010101111",  "000000010010100111",  "000000010010100000",  "000000010010011000",  "000000010010010001",  "000000010010001010",  "000000010010000010",  "000000010001111011",  "000000010001110011",  "000000010001101100",  "000000010001100100",  "000000010001011101",  "000000010001010101",  "000000010001001110",  "000000010001000110",  "000000010000111110",  "000000010000110111",  "000000010000101111",  "000000010000101000",  "000000010000100000",  "000000010000011000",  "000000010000010001",  "000000010000001001",  "000000010000000001",  "000000001111111010",  "000000001111110010",  "000000001111101010",  "000000001111100010",  "000000001111011011",  "000000001111010011",  "000000001111001011",  "000000001111000011",  "000000001110111100",  "000000001110110100",  "000000001110101100",  "000000001110100100",  "000000001110011100",  "000000001110010101",  "000000001110001101",  "000000001110000101",  "000000001101111101",  "000000001101110101",  "000000001101101101",  "000000001101100101",  "000000001101011101",  "000000001101010101",  "000000001101001101",  "000000001101000101",  "000000001100111101",  "000000001100110101",  "000000001100101110",  "000000001100100110",  "000000001100011101",  "000000001100010101",  "000000001100001101",  "000000001100000101",  "000000001011111101",  "000000001011110101",  "000000001011101101",  "000000001011100101",  "000000001011011101",  "000000001011010101",  "000000001011001101",  "000000001011000101",  "000000001010111101",  "000000001010110100",  "000000001010101100",  "000000001010100100",  "000000001010011100",  "000000001010010100",  "000000001010001100",  "000000001010000011",  "000000001001111011",  "000000001001110011",  "000000001001101011",  "000000001001100011",  "000000001001011010",  "000000001001010010",  "000000001001001010",  "000000001001000010",  "000000001000111001",  "000000001000110001",  "000000001000101001",  "000000001000100000",  "000000001000011000",  "000000001000010000",  "000000001000000111",  "000000000111111111",  "000000000111110111",  "000000000111101110",  "000000000111100110",  "000000000111011110",  "000000000111010101",  "000000000111001101",  "000000000111000101",  "000000000110111100",  "000000000110110100",  "000000000110101011",  "000000000110100011",  "000000000110011011",  "000000000110010010",  "000000000110001010",  "000000000110000001",  "000000000101111001",  "000000000101110000",  "000000000101101000",  "000000000101100000",  "000000000101010111",  "000000000101001111",  "000000000101000110",  "000000000100111110",  "000000000100110101",  "000000000100101101",  "000000000100100100",  "000000000100011100",  "000000000100010011",  "000000000100001011",  "000000000100000010",  "000000000011111001",  "000000000011110001",  "000000000011101000",  "000000000011100000",  "000000000011010111",  "000000000011001111",  "000000000011000110",  "000000000010111110",  "000000000010110101",  "000000000010101100",  "000000000010100100",  "000000000010011011",  "000000000010010011",  "000000000010001010",  "000000000010000001",  "000000000001111001",  "000000000001110000",  "000000000001101000",  "000000000001011111",  "000000000001010110",  "000000000001001110",  "000000000001000101",  "000000000000111101",  "000000000000110100",  "000000000000101011",  "000000000000100011",  "000000000000011010",  "000000000000010001",  "000000000000001001"),("000000000000000000",  "111111111111110111",  "111111111111101111",  "111111111111100110",  "111111111111011101",  "111111111111010101",  "111111111111001100",  "111111111111000011",  "111111111110111011",  "111111111110110010",  "111111111110101001",  "111111111110100001",  "111111111110011000",  "111111111110001111",  "111111111110000111",  "111111111101111110",  "111111111101110101",  "111111111101101100",  "111111111101100100",  "111111111101011011",  "111111111101010010",  "111111111101001010",  "111111111101000001",  "111111111100111000",  "111111111100110000",  "111111111100100111",  "111111111100011110",  "111111111100010101",  "111111111100001101",  "111111111100000100",  "111111111011111011",  "111111111011110011",  "111111111011101010",  "111111111011100001",  "111111111011011000",  "111111111011010000",  "111111111011000111",  "111111111010111110",  "111111111010110110",  "111111111010101101",  "111111111010100100",  "111111111010011011",  "111111111010010011",  "111111111010001010",  "111111111010000001",  "111111111001111001",  "111111111001110000",  "111111111001100111",  "111111111001011110",  "111111111001010110",  "111111111001001101",  "111111111001000100",  "111111111000111100",  "111111111000110011",  "111111111000101010",  "111111111000100001",  "111111111000011001",  "111111111000010000",  "111111111000000111",  "111111110111111111",  "111111110111110110",  "111111110111101101",  "111111110111100101",  "111111110111011100",  "111111110111010011",  "111111110111001010",  "111111110111000010",  "111111110110111001",  "111111110110110000",  "111111110110101000",  "111111110110011111",  "111111110110010110",  "111111110110001110",  "111111110110000101",  "111111110101111100",  "111111110101110100",  "111111110101101011",  "111111110101100010",  "111111110101011010",  "111111110101010001",  "111111110101001001",  "111111110101000000",  "111111110100110111",  "111111110100101111",  "111111110100100110",  "111111110100011101",  "111111110100010101",  "111111110100001100",  "111111110100000100",  "111111110011111011",  "111111110011110010",  "111111110011101010",  "111111110011100001",  "111111110011011001",  "111111110011010000",  "111111110011000111",  "111111110010111111",  "111111110010110110",  "111111110010101110",  "111111110010100101",  "111111110010011101",  "111111110010010100",  "111111110010001011",  "111111110010000011",  "111111110001111010",  "111111110001110010",  "111111110001101001",  "111111110001100001",  "111111110001011000",  "111111110001010000",  "111111110001000111",  "111111110000111111",  "111111110000110110",  "111111110000101110",  "111111110000100101",  "111111110000011101",  "111111110000010100",  "111111110000001100",  "111111110000000011",  "111111101111111011",  "111111101111110011",  "111111101111101010",  "111111101111100010",  "111111101111011001",  "111111101111010001",  "111111101111001001",  "111111101111000000",  "111111101110111000",  "111111101110101111",  "111111101110100111",  "111111101110011111",  "111111101110010110",  "111111101110001110",  "111111101110000110",  "111111101101111101",  "111111101101110101",  "111111101101101101",  "111111101101100100",  "111111101101011100",  "111111101101010100",  "111111101101001011",  "111111101101000011",  "111111101100111011",  "111111101100110011",  "111111101100101010",  "111111101100100010",  "111111101100011010",  "111111101100010010",  "111111101100001001",  "111111101100000001",  "111111101011111001",  "111111101011110001",  "111111101011101001",  "111111101011100000",  "111111101011011000",  "111111101011010000",  "111111101011001000",  "111111101011000000",  "111111101010111000",  "111111101010110000",  "111111101010101000",  "111111101010011111",  "111111101010010111",  "111111101010001111",  "111111101010000111",  "111111101001111111",  "111111101001110111",  "111111101001101111",  "111111101001100111",  "111111101001011111",  "111111101001010111",  "111111101001001111",  "111111101001000111",  "111111101000111111",  "111111101000110111",  "111111101000101111",  "111111101000100111",  "111111101000011111",  "111111101000011000",  "111111101000010000",  "111111101000001000",  "111111101000000000",  "111111100111111000",  "111111100111110000",  "111111100111101000",  "111111100111100001",  "111111100111011001",  "111111100111010001",  "111111100111001001",  "111111100111000001",  "111111100110111010",  "111111100110110010",  "111111100110101010",  "111111100110100010",  "111111100110011011",  "111111100110010011",  "111111100110001011",  "111111100110000100",  "111111100101111100",  "111111100101110100",  "111111100101101101",  "111111100101100101",  "111111100101011101",  "111111100101010110",  "111111100101001110",  "111111100101000111",  "111111100100111111",  "111111100100111000",  "111111100100110000",  "111111100100101000",  "111111100100100001",  "111111100100011010",  "111111100100010010",  "111111100100001011",  "111111100100000011",  "111111100011111100",  "111111100011110100",  "111111100011101101",  "111111100011100101",  "111111100011011110",  "111111100011010111",  "111111100011001111",  "111111100011001000",  "111111100011000001",  "111111100010111001",  "111111100010110010",  "111111100010101011",  "111111100010100100",  "111111100010011100",  "111111100010010101",  "111111100010001110",  "111111100010000111",  "111111100010000000",  "111111100001111000",  "111111100001110001",  "111111100001101010",  "111111100001100011",  "111111100001011100",  "111111100001010101",  "111111100001001110",  "111111100001000111",  "111111100001000000",  "111111100000111001",  "111111100000110010",  "111111100000101011",  "111111100000100100",  "111111100000011101",  "111111100000010110",  "111111100000001111",  "111111100000001000",  "111111100000000001",  "111111011111111010",  "111111011111110011",  "111111011111101101",  "111111011111100110",  "111111011111011111",  "111111011111011000",  "111111011111010001",  "111111011111001011",  "111111011111000100",  "111111011110111101",  "111111011110110111",  "111111011110110000",  "111111011110101001",  "111111011110100011",  "111111011110011100",  "111111011110010101",  "111111011110001111",  "111111011110001000",  "111111011110000010",  "111111011101111011",  "111111011101110101",  "111111011101101110",  "111111011101101000",  "111111011101100001",  "111111011101011011",  "111111011101010100",  "111111011101001110",  "111111011101001000",  "111111011101000001",  "111111011100111011",  "111111011100110100",  "111111011100101110",  "111111011100101000",  "111111011100100010",  "111111011100011011",  "111111011100010101",  "111111011100001111",  "111111011100001001",  "111111011100000011",  "111111011011111100",  "111111011011110110",  "111111011011110000",  "111111011011101010",  "111111011011100100",  "111111011011011110",  "111111011011011000",  "111111011011010010",  "111111011011001100",  "111111011011000110",  "111111011011000000",  "111111011010111010",  "111111011010110100",  "111111011010101110",  "111111011010101000",  "111111011010100010",  "111111011010011101",  "111111011010010111",  "111111011010010001",  "111111011010001011",  "111111011010000101",  "111111011010000000",  "111111011001111010",  "111111011001110100",  "111111011001101111",  "111111011001101001",  "111111011001100011",  "111111011001011110",  "111111011001011000",  "111111011001010011",  "111111011001001101",  "111111011001001000",  "111111011001000010",  "111111011000111101",  "111111011000110111",  "111111011000110010",  "111111011000101100",  "111111011000100111",  "111111011000100010",  "111111011000011100",  "111111011000010111",  "111111011000010010",  "111111011000001100",  "111111011000000111",  "111111011000000010",  "111111010111111101",  "111111010111110111",  "111111010111110010",  "111111010111101101",  "111111010111101000",  "111111010111100011",  "111111010111011110",  "111111010111011001",  "111111010111010100",  "111111010111001111",  "111111010111001010",  "111111010111000101",  "111111010111000000",  "111111010110111011",  "111111010110110110",  "111111010110110001",  "111111010110101100",  "111111010110101000",  "111111010110100011",  "111111010110011110",  "111111010110011001",  "111111010110010101",  "111111010110010000",  "111111010110001011",  "111111010110000110",  "111111010110000010",  "111111010101111101",  "111111010101111001",  "111111010101110100",  "111111010101110000",  "111111010101101011",  "111111010101100111",  "111111010101100010",  "111111010101011110",  "111111010101011001",  "111111010101010101",  "111111010101010000",  "111111010101001100",  "111111010101001000",  "111111010101000011",  "111111010100111111",  "111111010100111011",  "111111010100110111",  "111111010100110011",  "111111010100101110",  "111111010100101010",  "111111010100100110",  "111111010100100010",  "111111010100011110",  "111111010100011010",  "111111010100010110",  "111111010100010010",  "111111010100001110",  "111111010100001010",  "111111010100000110",  "111111010100000010",  "111111010011111110",  "111111010011111010",  "111111010011110110",  "111111010011110011",  "111111010011101111",  "111111010011101011",  "111111010011100111",  "111111010011100100",  "111111010011100000",  "111111010011011100",  "111111010011011001",  "111111010011010101",  "111111010011010010",  "111111010011001110",  "111111010011001011",  "111111010011000111",  "111111010011000100",  "111111010011000000",  "111111010010111101",  "111111010010111001",  "111111010010110110",  "111111010010110011",  "111111010010101111",  "111111010010101100",  "111111010010101001",  "111111010010100110",  "111111010010100010",  "111111010010011111",  "111111010010011100",  "111111010010011001",  "111111010010010110",  "111111010010010011",  "111111010010010000",  "111111010010001101",  "111111010010001010",  "111111010010000111",  "111111010010000100",  "111111010010000001",  "111111010001111110",  "111111010001111011",  "111111010001111000",  "111111010001110101",  "111111010001110011",  "111111010001110000",  "111111010001101101",  "111111010001101011",  "111111010001101000",  "111111010001100101",  "111111010001100011",  "111111010001100000",  "111111010001011101",  "111111010001011011",  "111111010001011000",  "111111010001010110",  "111111010001010011",  "111111010001010001",  "111111010001001111",  "111111010001001100",  "111111010001001010",  "111111010001001000",  "111111010001000101",  "111111010001000011",  "111111010001000001",  "111111010000111111",  "111111010000111100",  "111111010000111010",  "111111010000111000",  "111111010000110110",  "111111010000110100",  "111111010000110010",  "111111010000110000",  "111111010000101110",  "111111010000101100",  "111111010000101010",  "111111010000101000",  "111111010000100110",  "111111010000100100",  "111111010000100011",  "111111010000100001",  "111111010000011111",  "111111010000011101",  "111111010000011100",  "111111010000011010",  "111111010000011000",  "111111010000010111",  "111111010000010101",  "111111010000010100",  "111111010000010010",  "111111010000010000",  "111111010000001111",  "111111010000001110",  "111111010000001100",  "111111010000001011",  "111111010000001001",  "111111010000001000",  "111111010000000111",  "111111010000000101",  "111111010000000100",  "111111010000000011",  "111111010000000010",  "111111010000000001",  "111111001111111111",  "111111001111111110",  "111111001111111101",  "111111001111111100",  "111111001111111011",  "111111001111111010",  "111111001111111001",  "111111001111111000",  "111111001111110111",  "111111001111110111",  "111111001111110110",  "111111001111110101",  "111111001111110100",  "111111001111110011",  "111111001111110011",  "111111001111110010",  "111111001111110001",  "111111001111110001",  "111111001111110000",  "111111001111101111",  "111111001111101111",  "111111001111101110",  "111111001111101110",  "111111001111101101",  "111111001111101101",  "111111001111101100",  "111111001111101100",  "111111001111101100",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101100",  "111111001111101100",  "111111001111101101",  "111111001111101101",  "111111001111101101",  "111111001111101110",  "111111001111101110",  "111111001111101111",  "111111001111110000",  "111111001111110000",  "111111001111110001",  "111111001111110010",  "111111001111110010",  "111111001111110011",  "111111001111110100",  "111111001111110100",  "111111001111110101",  "111111001111110110",  "111111001111110111",  "111111001111111000",  "111111001111111001",  "111111001111111010",  "111111001111111011",  "111111001111111100",  "111111001111111101",  "111111001111111110",  "111111001111111111",  "111111010000000000",  "111111010000000001",  "111111010000000011",  "111111010000000100",  "111111010000000101",  "111111010000000110",  "111111010000001000",  "111111010000001001",  "111111010000001010",  "111111010000001100",  "111111010000001101",  "111111010000001111",  "111111010000010000",  "111111010000010010",  "111111010000010011",  "111111010000010101",  "111111010000010110",  "111111010000011000",  "111111010000011010",  "111111010000011011",  "111111010000011101",  "111111010000011111",  "111111010000100001",  "111111010000100010",  "111111010000100100",  "111111010000100110",  "111111010000101000",  "111111010000101010",  "111111010000101100",  "111111010000101110",  "111111010000110000",  "111111010000110010",  "111111010000110100",  "111111010000110110",  "111111010000111000",  "111111010000111010",  "111111010000111101",  "111111010000111111",  "111111010001000001",  "111111010001000011",  "111111010001000110",  "111111010001001000",  "111111010001001010",  "111111010001001101",  "111111010001001111",  "111111010001010010",  "111111010001010100",  "111111010001010111",  "111111010001011001",  "111111010001011100",  "111111010001011110",  "111111010001100001",  "111111010001100100",  "111111010001100110",  "111111010001101001",  "111111010001101100",  "111111010001101111",  "111111010001110001",  "111111010001110100",  "111111010001110111",  "111111010001111010",  "111111010001111101",  "111111010010000000",  "111111010010000011",  "111111010010000110",  "111111010010001001",  "111111010010001100",  "111111010010001111",  "111111010010010010",  "111111010010010101",  "111111010010011000",  "111111010010011100",  "111111010010011111",  "111111010010100010",  "111111010010100101",  "111111010010101001",  "111111010010101100",  "111111010010110000",  "111111010010110011",  "111111010010110110",  "111111010010111010",  "111111010010111101",  "111111010011000001",  "111111010011000100",  "111111010011001000",  "111111010011001100",  "111111010011001111",  "111111010011010011",  "111111010011010111",  "111111010011011010",  "111111010011011110",  "111111010011100010",  "111111010011100110",  "111111010011101001",  "111111010011101101",  "111111010011110001",  "111111010011110101",  "111111010011111001",  "111111010011111101",  "111111010100000001",  "111111010100000101",  "111111010100001001",  "111111010100001101",  "111111010100010001",  "111111010100010101",  "111111010100011010",  "111111010100011110",  "111111010100100010",  "111111010100100110",  "111111010100101011",  "111111010100101111",  "111111010100110011",  "111111010100111000",  "111111010100111100",  "111111010101000000",  "111111010101000101",  "111111010101001001",  "111111010101001110",  "111111010101010010",  "111111010101010111",  "111111010101011011",  "111111010101100000",  "111111010101100101",  "111111010101101001",  "111111010101101110",  "111111010101110011",  "111111010101111000",  "111111010101111100",  "111111010110000001",  "111111010110000110",  "111111010110001011",  "111111010110010000",  "111111010110010101",  "111111010110011010",  "111111010110011110",  "111111010110100011",  "111111010110101000",  "111111010110101110",  "111111010110110011",  "111111010110111000",  "111111010110111101",  "111111010111000010",  "111111010111000111",  "111111010111001100",  "111111010111010010",  "111111010111010111",  "111111010111011100",  "111111010111100001",  "111111010111100111",  "111111010111101100",  "111111010111110010",  "111111010111110111",  "111111010111111100",  "111111011000000010",  "111111011000000111",  "111111011000001101",  "111111011000010010",  "111111011000011000",  "111111011000011110",  "111111011000100011",  "111111011000101001",  "111111011000101110",  "111111011000110100",  "111111011000111010",  "111111011001000000",  "111111011001000101",  "111111011001001011",  "111111011001010001",  "111111011001010111",  "111111011001011101",  "111111011001100011",  "111111011001101001",  "111111011001101111",  "111111011001110101",  "111111011001111011",  "111111011010000001",  "111111011010000111",  "111111011010001101",  "111111011010010011",  "111111011010011001",  "111111011010011111",  "111111011010100101",  "111111011010101100",  "111111011010110010",  "111111011010111000",  "111111011010111110",  "111111011011000101",  "111111011011001011",  "111111011011010001",  "111111011011011000",  "111111011011011110",  "111111011011100100",  "111111011011101011",  "111111011011110001",  "111111011011111000",  "111111011011111110",  "111111011100000101",  "111111011100001100",  "111111011100010010",  "111111011100011001",  "111111011100011111",  "111111011100100110",  "111111011100101101",  "111111011100110011",  "111111011100111010",  "111111011101000001",  "111111011101001000",  "111111011101001111",  "111111011101010101",  "111111011101011100",  "111111011101100011",  "111111011101101010",  "111111011101110001",  "111111011101111000",  "111111011101111111",  "111111011110000110",  "111111011110001101",  "111111011110010100",  "111111011110011011",  "111111011110100010",  "111111011110101001",  "111111011110110000",  "111111011110110111",  "111111011110111111",  "111111011111000110",  "111111011111001101",  "111111011111010100",  "111111011111011100",  "111111011111100011",  "111111011111101010",  "111111011111110001",  "111111011111111001",  "111111100000000000",  "111111100000001000",  "111111100000001111",  "111111100000010110",  "111111100000011110",  "111111100000100101",  "111111100000101101",  "111111100000110100",  "111111100000111100",  "111111100001000100",  "111111100001001011",  "111111100001010011",  "111111100001011010",  "111111100001100010",  "111111100001101010",  "111111100001110001",  "111111100001111001",  "111111100010000001",  "111111100010001001",  "111111100010010000",  "111111100010011000",  "111111100010100000",  "111111100010101000",  "111111100010110000",  "111111100010111000",  "111111100011000000",  "111111100011001000",  "111111100011001111",  "111111100011010111",  "111111100011011111",  "111111100011100111",  "111111100011101111",  "111111100011111000",  "111111100100000000",  "111111100100001000",  "111111100100010000",  "111111100100011000",  "111111100100100000",  "111111100100101000",  "111111100100110000",  "111111100100111001",  "111111100101000001",  "111111100101001001",  "111111100101010001",  "111111100101011010",  "111111100101100010",  "111111100101101010",  "111111100101110011",  "111111100101111011",  "111111100110000011",  "111111100110001100",  "111111100110010100",  "111111100110011101",  "111111100110100101",  "111111100110101101",  "111111100110110110",  "111111100110111110",  "111111100111000111",  "111111100111010000",  "111111100111011000",  "111111100111100001",  "111111100111101001",  "111111100111110010",  "111111100111111011",  "111111101000000011",  "111111101000001100",  "111111101000010101",  "111111101000011101",  "111111101000100110",  "111111101000101111",  "111111101000110111",  "111111101001000000",  "111111101001001001",  "111111101001010010",  "111111101001011011",  "111111101001100011",  "111111101001101100",  "111111101001110101",  "111111101001111110",  "111111101010000111",  "111111101010010000",  "111111101010011001",  "111111101010100010",  "111111101010101011",  "111111101010110100",  "111111101010111101",  "111111101011000110",  "111111101011001111",  "111111101011011000",  "111111101011100001",  "111111101011101010",  "111111101011110011",  "111111101011111100",  "111111101100000101",  "111111101100001110",  "111111101100011000",  "111111101100100001",  "111111101100101010",  "111111101100110011",  "111111101100111100",  "111111101101000110",  "111111101101001111",  "111111101101011000",  "111111101101100001",  "111111101101101011",  "111111101101110100",  "111111101101111101",  "111111101110000111",  "111111101110010000",  "111111101110011001",  "111111101110100011",  "111111101110101100",  "111111101110110101",  "111111101110111111",  "111111101111001000",  "111111101111010010",  "111111101111011011",  "111111101111100101",  "111111101111101110",  "111111101111111000",  "111111110000000001",  "111111110000001011",  "111111110000010100",  "111111110000011110",  "111111110000100111",  "111111110000110001",  "111111110000111010",  "111111110001000100",  "111111110001001110",  "111111110001010111",  "111111110001100001",  "111111110001101011",  "111111110001110100",  "111111110001111110",  "111111110010001000",  "111111110010010001",  "111111110010011011",  "111111110010100101",  "111111110010101110",  "111111110010111000",  "111111110011000010",  "111111110011001100",  "111111110011010110",  "111111110011011111",  "111111110011101001",  "111111110011110011",  "111111110011111101",  "111111110100000111",  "111111110100010000",  "111111110100011010",  "111111110100100100",  "111111110100101110",  "111111110100111000",  "111111110101000010",  "111111110101001100",  "111111110101010110",  "111111110101100000",  "111111110101101001",  "111111110101110011",  "111111110101111101",  "111111110110000111",  "111111110110010001",  "111111110110011011",  "111111110110100101",  "111111110110101111",  "111111110110111001",  "111111110111000011",  "111111110111001101",  "111111110111010111",  "111111110111100001",  "111111110111101011",  "111111110111110110",  "111111111000000000",  "111111111000001010",  "111111111000010100",  "111111111000011110",  "111111111000101000",  "111111111000110010",  "111111111000111100",  "111111111001000110",  "111111111001010000",  "111111111001011011",  "111111111001100101",  "111111111001101111",  "111111111001111001",  "111111111010000011",  "111111111010001101",  "111111111010011000",  "111111111010100010",  "111111111010101100",  "111111111010110110",  "111111111011000000",  "111111111011001011",  "111111111011010101",  "111111111011011111",  "111111111011101001",  "111111111011110100",  "111111111011111110",  "111111111100001000",  "111111111100010010",  "111111111100011101",  "111111111100100111",  "111111111100110001",  "111111111100111100",  "111111111101000110",  "111111111101010000",  "111111111101011010",  "111111111101100101",  "111111111101101111",  "111111111101111001",  "111111111110000100",  "111111111110001110",  "111111111110011000",  "111111111110100011",  "111111111110101101",  "111111111110110111",  "111111111111000010",  "111111111111001100",  "111111111111010111",  "111111111111100001",  "111111111111101011",  "111111111111110110"),("000000000000000000",  "000000000000001010",  "000000000000010101",  "000000000000011111",  "000000000000101010",  "000000000000110100",  "000000000000111110",  "000000000001001001",  "000000000001010011",  "000000000001011110",  "000000000001101000",  "000000000001110010",  "000000000001111101",  "000000000010000111",  "000000000010010010",  "000000000010011100",  "000000000010100110",  "000000000010110001",  "000000000010111011",  "000000000011000110",  "000000000011010000",  "000000000011011011",  "000000000011100101",  "000000000011110000",  "000000000011111010",  "000000000100000100",  "000000000100001111",  "000000000100011001",  "000000000100100100",  "000000000100101110",  "000000000100111001",  "000000000101000011",  "000000000101001110",  "000000000101011000",  "000000000101100010",  "000000000101101101",  "000000000101110111",  "000000000110000010",  "000000000110001100",  "000000000110010111",  "000000000110100001",  "000000000110101100",  "000000000110110110",  "000000000111000000",  "000000000111001011",  "000000000111010101",  "000000000111100000",  "000000000111101010",  "000000000111110101",  "000000000111111111",  "000000001000001010",  "000000001000010100",  "000000001000011111",  "000000001000101001",  "000000001000110011",  "000000001000111110",  "000000001001001000",  "000000001001010011",  "000000001001011101",  "000000001001101000",  "000000001001110010",  "000000001001111100",  "000000001010000111",  "000000001010010001",  "000000001010011100",  "000000001010100110",  "000000001010110001",  "000000001010111011",  "000000001011000101",  "000000001011010000",  "000000001011011010",  "000000001011100101",  "000000001011101111",  "000000001011111001",  "000000001100000100",  "000000001100001110",  "000000001100011000",  "000000001100100011",  "000000001100101101",  "000000001100111000",  "000000001101000010",  "000000001101001100",  "000000001101010111",  "000000001101100001",  "000000001101101011",  "000000001101110110",  "000000001110000000",  "000000001110001010",  "000000001110010101",  "000000001110011111",  "000000001110101001",  "000000001110110100",  "000000001110111110",  "000000001111001000",  "000000001111010011",  "000000001111011101",  "000000001111100111",  "000000001111110001",  "000000001111111100",  "000000010000000110",  "000000010000010000",  "000000010000011011",  "000000010000100101",  "000000010000101111",  "000000010000111001",  "000000010001000011",  "000000010001001110",  "000000010001011000",  "000000010001100010",  "000000010001101100",  "000000010001110111",  "000000010010000001",  "000000010010001011",  "000000010010010101",  "000000010010011111",  "000000010010101001",  "000000010010110100",  "000000010010111110",  "000000010011001000",  "000000010011010010",  "000000010011011100",  "000000010011100110",  "000000010011110000",  "000000010011111010",  "000000010100000100",  "000000010100001111",  "000000010100011001",  "000000010100100011",  "000000010100101101",  "000000010100110111",  "000000010101000001",  "000000010101001011",  "000000010101010101",  "000000010101011111",  "000000010101101001",  "000000010101110011",  "000000010101111101",  "000000010110000111",  "000000010110010001",  "000000010110011011",  "000000010110100101",  "000000010110101111",  "000000010110111001",  "000000010111000010",  "000000010111001100",  "000000010111010110",  "000000010111100000",  "000000010111101010",  "000000010111110100",  "000000010111111110",  "000000011000001000",  "000000011000010001",  "000000011000011011",  "000000011000100101",  "000000011000101111",  "000000011000111001",  "000000011001000010",  "000000011001001100",  "000000011001010110",  "000000011001100000",  "000000011001101001",  "000000011001110011",  "000000011001111101",  "000000011010000110",  "000000011010010000",  "000000011010011010",  "000000011010100011",  "000000011010101101",  "000000011010110111",  "000000011011000000",  "000000011011001010",  "000000011011010011",  "000000011011011101",  "000000011011100110",  "000000011011110000",  "000000011011111010",  "000000011100000011",  "000000011100001101",  "000000011100010110",  "000000011100100000",  "000000011100101001",  "000000011100110010",  "000000011100111100",  "000000011101000101",  "000000011101001111",  "000000011101011000",  "000000011101100001",  "000000011101101011",  "000000011101110100",  "000000011101111110",  "000000011110000111",  "000000011110010000",  "000000011110011001",  "000000011110100011",  "000000011110101100",  "000000011110110101",  "000000011110111110",  "000000011111001000",  "000000011111010001",  "000000011111011010",  "000000011111100011",  "000000011111101100",  "000000011111110101",  "000000011111111111",  "000000100000001000",  "000000100000010001",  "000000100000011010",  "000000100000100011",  "000000100000101100",  "000000100000110101",  "000000100000111110",  "000000100001000111",  "000000100001010000",  "000000100001011001",  "000000100001100010",  "000000100001101011",  "000000100001110100",  "000000100001111101",  "000000100010000101",  "000000100010001110",  "000000100010010111",  "000000100010100000",  "000000100010101001",  "000000100010110001",  "000000100010111010",  "000000100011000011",  "000000100011001100",  "000000100011010100",  "000000100011011101",  "000000100011100110",  "000000100011101110",  "000000100011110111",  "000000100100000000",  "000000100100001000",  "000000100100010001",  "000000100100011001",  "000000100100100010",  "000000100100101010",  "000000100100110011",  "000000100100111011",  "000000100101000100",  "000000100101001100",  "000000100101010101",  "000000100101011101",  "000000100101100110",  "000000100101101110",  "000000100101110110",  "000000100101111111",  "000000100110000111",  "000000100110001111",  "000000100110010111",  "000000100110100000",  "000000100110101000",  "000000100110110000",  "000000100110111000",  "000000100111000001",  "000000100111001001",  "000000100111010001",  "000000100111011001",  "000000100111100001",  "000000100111101001",  "000000100111110001",  "000000100111111001",  "000000101000000001",  "000000101000001001",  "000000101000010001",  "000000101000011001",  "000000101000100001",  "000000101000101001",  "000000101000110001",  "000000101000111000",  "000000101001000000",  "000000101001001000",  "000000101001010000",  "000000101001011000",  "000000101001011111",  "000000101001100111",  "000000101001101111",  "000000101001110110",  "000000101001111110",  "000000101010000110",  "000000101010001101",  "000000101010010101",  "000000101010011100",  "000000101010100100",  "000000101010101011",  "000000101010110011",  "000000101010111010",  "000000101011000010",  "000000101011001001",  "000000101011010001",  "000000101011011000",  "000000101011011111",  "000000101011100111",  "000000101011101110",  "000000101011110101",  "000000101011111101",  "000000101100000100",  "000000101100001011",  "000000101100010010",  "000000101100011001",  "000000101100100000",  "000000101100101000",  "000000101100101111",  "000000101100110110",  "000000101100111101",  "000000101101000100",  "000000101101001011",  "000000101101010010",  "000000101101011001",  "000000101101100000",  "000000101101100110",  "000000101101101101",  "000000101101110100",  "000000101101111011",  "000000101110000010",  "000000101110001000",  "000000101110001111",  "000000101110010110",  "000000101110011101",  "000000101110100011",  "000000101110101010",  "000000101110110000",  "000000101110110111",  "000000101110111110",  "000000101111000100",  "000000101111001011",  "000000101111010001",  "000000101111011000",  "000000101111011110",  "000000101111100100",  "000000101111101011",  "000000101111110001",  "000000101111110111",  "000000101111111110",  "000000110000000100",  "000000110000001010",  "000000110000010000",  "000000110000010111",  "000000110000011101",  "000000110000100011",  "000000110000101001",  "000000110000101111",  "000000110000110101",  "000000110000111011",  "000000110001000001",  "000000110001000111",  "000000110001001101",  "000000110001010011",  "000000110001011001",  "000000110001011111",  "000000110001100100",  "000000110001101010",  "000000110001110000",  "000000110001110110",  "000000110001111011",  "000000110010000001",  "000000110010000111",  "000000110010001100",  "000000110010010010",  "000000110010011000",  "000000110010011101",  "000000110010100011",  "000000110010101000",  "000000110010101110",  "000000110010110011",  "000000110010111000",  "000000110010111110",  "000000110011000011",  "000000110011001000",  "000000110011001110",  "000000110011010011",  "000000110011011000",  "000000110011011101",  "000000110011100011",  "000000110011101000",  "000000110011101101",  "000000110011110010",  "000000110011110111",  "000000110011111100",  "000000110100000001",  "000000110100000110",  "000000110100001011",  "000000110100010000",  "000000110100010101",  "000000110100011010",  "000000110100011110",  "000000110100100011",  "000000110100101000",  "000000110100101101",  "000000110100110001",  "000000110100110110",  "000000110100111011",  "000000110100111111",  "000000110101000100",  "000000110101001000",  "000000110101001101",  "000000110101010001",  "000000110101010110",  "000000110101011010",  "000000110101011111",  "000000110101100011",  "000000110101100111",  "000000110101101100",  "000000110101110000",  "000000110101110100",  "000000110101111000",  "000000110101111100",  "000000110110000001",  "000000110110000101",  "000000110110001001",  "000000110110001101",  "000000110110010001",  "000000110110010101",  "000000110110011001",  "000000110110011101",  "000000110110100001",  "000000110110100100",  "000000110110101000",  "000000110110101100",  "000000110110110000",  "000000110110110100",  "000000110110110111",  "000000110110111011",  "000000110110111111",  "000000110111000010",  "000000110111000110",  "000000110111001001",  "000000110111001101",  "000000110111010000",  "000000110111010100",  "000000110111010111",  "000000110111011010",  "000000110111011110",  "000000110111100001",  "000000110111100100",  "000000110111101000",  "000000110111101011",  "000000110111101110",  "000000110111110001",  "000000110111110100",  "000000110111110111",  "000000110111111011",  "000000110111111110",  "000000111000000001",  "000000111000000011",  "000000111000000110",  "000000111000001001",  "000000111000001100",  "000000111000001111",  "000000111000010010",  "000000111000010101",  "000000111000010111",  "000000111000011010",  "000000111000011101",  "000000111000011111",  "000000111000100010",  "000000111000100100",  "000000111000100111",  "000000111000101001",  "000000111000101100",  "000000111000101110",  "000000111000110001",  "000000111000110011",  "000000111000110101",  "000000111000111000",  "000000111000111010",  "000000111000111100",  "000000111000111110",  "000000111001000001",  "000000111001000011",  "000000111001000101",  "000000111001000111",  "000000111001001001",  "000000111001001011",  "000000111001001101",  "000000111001001111",  "000000111001010001",  "000000111001010010",  "000000111001010100",  "000000111001010110",  "000000111001011000",  "000000111001011010",  "000000111001011011",  "000000111001011101",  "000000111001011111",  "000000111001100000",  "000000111001100010",  "000000111001100011",  "000000111001100101",  "000000111001100110",  "000000111001101000",  "000000111001101001",  "000000111001101010",  "000000111001101100",  "000000111001101101",  "000000111001101110",  "000000111001101111",  "000000111001110000",  "000000111001110010",  "000000111001110011",  "000000111001110100",  "000000111001110101",  "000000111001110110",  "000000111001110111",  "000000111001111000",  "000000111001111001",  "000000111001111001",  "000000111001111010",  "000000111001111011",  "000000111001111100",  "000000111001111101",  "000000111001111101",  "000000111001111110",  "000000111001111110",  "000000111001111111",  "000000111010000000",  "000000111010000000",  "000000111010000001",  "000000111010000001",  "000000111010000001",  "000000111010000010",  "000000111010000010",  "000000111010000010",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000010",  "000000111010000010",  "000000111010000010",  "000000111010000001",  "000000111010000001",  "000000111010000000",  "000000111010000000",  "000000111001111111",  "000000111001111111",  "000000111001111110",  "000000111001111101",  "000000111001111101",  "000000111001111100",  "000000111001111011",  "000000111001111011",  "000000111001111010",  "000000111001111001",  "000000111001111000",  "000000111001110111",  "000000111001110110",  "000000111001110101",  "000000111001110100",  "000000111001110011",  "000000111001110010",  "000000111001110001",  "000000111001110000",  "000000111001101110",  "000000111001101101",  "000000111001101100",  "000000111001101010",  "000000111001101001",  "000000111001101000",  "000000111001100110",  "000000111001100101",  "000000111001100011",  "000000111001100010",  "000000111001100000",  "000000111001011111",  "000000111001011101",  "000000111001011011",  "000000111001011010",  "000000111001011000",  "000000111001010110",  "000000111001010100",  "000000111001010011",  "000000111001010001",  "000000111001001111",  "000000111001001101",  "000000111001001011",  "000000111001001001",  "000000111001000111",  "000000111001000101",  "000000111001000011",  "000000111001000000",  "000000111000111110",  "000000111000111100",  "000000111000111010",  "000000111000110111",  "000000111000110101",  "000000111000110011",  "000000111000110000",  "000000111000101110",  "000000111000101011",  "000000111000101001",  "000000111000100110",  "000000111000100100",  "000000111000100001",  "000000111000011110",  "000000111000011100",  "000000111000011001",  "000000111000010110",  "000000111000010011",  "000000111000010001",  "000000111000001110",  "000000111000001011",  "000000111000001000",  "000000111000000101",  "000000111000000010",  "000000110111111111",  "000000110111111100",  "000000110111111001",  "000000110111110110",  "000000110111110010",  "000000110111101111",  "000000110111101100",  "000000110111101001",  "000000110111100101",  "000000110111100010",  "000000110111011111",  "000000110111011011",  "000000110111011000",  "000000110111010100",  "000000110111010001",  "000000110111001101",  "000000110111001001",  "000000110111000110",  "000000110111000010",  "000000110110111111",  "000000110110111011",  "000000110110110111",  "000000110110110011",  "000000110110101111",  "000000110110101011",  "000000110110101000",  "000000110110100100",  "000000110110100000",  "000000110110011100",  "000000110110011000",  "000000110110010100",  "000000110110001111",  "000000110110001011",  "000000110110000111",  "000000110110000011",  "000000110101111111",  "000000110101111010",  "000000110101110110",  "000000110101110010",  "000000110101101101",  "000000110101101001",  "000000110101100100",  "000000110101100000",  "000000110101011011",  "000000110101010111",  "000000110101010010",  "000000110101001110",  "000000110101001001",  "000000110101000100",  "000000110101000000",  "000000110100111011",  "000000110100110110",  "000000110100110001",  "000000110100101100",  "000000110100100111",  "000000110100100010",  "000000110100011110",  "000000110100011001",  "000000110100010011",  "000000110100001110",  "000000110100001001",  "000000110100000100",  "000000110011111111",  "000000110011111010",  "000000110011110101",  "000000110011101111",  "000000110011101010",  "000000110011100101",  "000000110011011111",  "000000110011011010",  "000000110011010101",  "000000110011001111",  "000000110011001010",  "000000110011000100",  "000000110010111111",  "000000110010111001",  "000000110010110011",  "000000110010101110",  "000000110010101000",  "000000110010100010",  "000000110010011100",  "000000110010010111",  "000000110010010001",  "000000110010001011",  "000000110010000101",  "000000110001111111",  "000000110001111001",  "000000110001110011",  "000000110001101101",  "000000110001100111",  "000000110001100001",  "000000110001011011",  "000000110001010101",  "000000110001001111",  "000000110001001001",  "000000110001000010",  "000000110000111100",  "000000110000110110",  "000000110000101111",  "000000110000101001",  "000000110000100011",  "000000110000011100",  "000000110000010110",  "000000110000001111",  "000000110000001001",  "000000110000000010",  "000000101111111100",  "000000101111110101",  "000000101111101110",  "000000101111101000",  "000000101111100001",  "000000101111011010",  "000000101111010011",  "000000101111001101",  "000000101111000110",  "000000101110111111",  "000000101110111000",  "000000101110110001",  "000000101110101010",  "000000101110100011",  "000000101110011100",  "000000101110010101",  "000000101110001110",  "000000101110000111",  "000000101110000000",  "000000101101111001",  "000000101101110001",  "000000101101101010",  "000000101101100011",  "000000101101011100",  "000000101101010100",  "000000101101001101",  "000000101101000101",  "000000101100111110",  "000000101100110111",  "000000101100101111",  "000000101100101000",  "000000101100100000",  "000000101100011001",  "000000101100010001",  "000000101100001001",  "000000101100000010",  "000000101011111010",  "000000101011110010",  "000000101011101011",  "000000101011100011",  "000000101011011011",  "000000101011010011",  "000000101011001011",  "000000101011000011",  "000000101010111011",  "000000101010110100",  "000000101010101100",  "000000101010100100",  "000000101010011100",  "000000101010010011",  "000000101010001011",  "000000101010000011",  "000000101001111011",  "000000101001110011",  "000000101001101011",  "000000101001100011",  "000000101001011010",  "000000101001010010",  "000000101001001010",  "000000101001000001",  "000000101000111001",  "000000101000110001",  "000000101000101000",  "000000101000100000",  "000000101000010111",  "000000101000001111",  "000000101000000110",  "000000100111111110",  "000000100111110101",  "000000100111101100",  "000000100111100100",  "000000100111011011",  "000000100111010010",  "000000100111001010",  "000000100111000001",  "000000100110111000",  "000000100110101111",  "000000100110100111",  "000000100110011110",  "000000100110010101",  "000000100110001100",  "000000100110000011",  "000000100101111010",  "000000100101110001",  "000000100101101000",  "000000100101011111",  "000000100101010110",  "000000100101001101",  "000000100101000100",  "000000100100111011",  "000000100100110001",  "000000100100101000",  "000000100100011111",  "000000100100010110",  "000000100100001100",  "000000100100000011",  "000000100011111010",  "000000100011110000",  "000000100011100111",  "000000100011011110",  "000000100011010100",  "000000100011001011",  "000000100011000001",  "000000100010111000",  "000000100010101110",  "000000100010100101",  "000000100010011011",  "000000100010010010",  "000000100010001000",  "000000100001111110",  "000000100001110101",  "000000100001101011",  "000000100001100001",  "000000100001011000",  "000000100001001110",  "000000100001000100",  "000000100000111010",  "000000100000110000",  "000000100000100111",  "000000100000011101",  "000000100000010011",  "000000100000001001",  "000000011111111111",  "000000011111110101",  "000000011111101011",  "000000011111100001",  "000000011111010111",  "000000011111001101",  "000000011111000011",  "000000011110111001",  "000000011110101110",  "000000011110100100",  "000000011110011010",  "000000011110010000",  "000000011110000110",  "000000011101111011",  "000000011101110001",  "000000011101100111",  "000000011101011101",  "000000011101010010",  "000000011101001000",  "000000011100111110",  "000000011100110011",  "000000011100101001",  "000000011100011110",  "000000011100010100",  "000000011100001001",  "000000011011111111",  "000000011011110100",  "000000011011101010",  "000000011011011111",  "000000011011010101",  "000000011011001010",  "000000011011000000",  "000000011010110101",  "000000011010101010",  "000000011010100000",  "000000011010010101",  "000000011010001010",  "000000011001111111",  "000000011001110101",  "000000011001101010",  "000000011001011111",  "000000011001010100",  "000000011001001001",  "000000011000111111",  "000000011000110100",  "000000011000101001",  "000000011000011110",  "000000011000010011",  "000000011000001000",  "000000010111111101",  "000000010111110010",  "000000010111100111",  "000000010111011100",  "000000010111010001",  "000000010111000110",  "000000010110111011",  "000000010110110000",  "000000010110100101",  "000000010110011010",  "000000010110001110",  "000000010110000011",  "000000010101111000",  "000000010101101101",  "000000010101100010",  "000000010101010110",  "000000010101001011",  "000000010101000000",  "000000010100110101",  "000000010100101001",  "000000010100011110",  "000000010100010011",  "000000010100000111",  "000000010011111100",  "000000010011110000",  "000000010011100101",  "000000010011011010",  "000000010011001110",  "000000010011000011",  "000000010010110111",  "000000010010101100",  "000000010010100000",  "000000010010010101",  "000000010010001001",  "000000010001111110",  "000000010001110010",  "000000010001100111",  "000000010001011011",  "000000010001001111",  "000000010001000100",  "000000010000111000",  "000000010000101101",  "000000010000100001",  "000000010000010101",  "000000010000001010",  "000000001111111110",  "000000001111110010",  "000000001111100110",  "000000001111011011",  "000000001111001111",  "000000001111000011",  "000000001110110111",  "000000001110101100",  "000000001110100000",  "000000001110010100",  "000000001110001000",  "000000001101111100",  "000000001101110000",  "000000001101100101",  "000000001101011001",  "000000001101001101",  "000000001101000001",  "000000001100110101",  "000000001100101001",  "000000001100011101",  "000000001100010001",  "000000001100000101",  "000000001011111001",  "000000001011101101",  "000000001011100001",  "000000001011010101",  "000000001011001001",  "000000001010111101",  "000000001010110001",  "000000001010100101",  "000000001010011001",  "000000001010001101",  "000000001010000001",  "000000001001110101",  "000000001001101000",  "000000001001011100",  "000000001001010000",  "000000001001000100",  "000000001000111000",  "000000001000101100",  "000000001000100000",  "000000001000010011",  "000000001000000111",  "000000000111111011",  "000000000111101111",  "000000000111100011",  "000000000111010110",  "000000000111001010",  "000000000110111110",  "000000000110110010",  "000000000110100101",  "000000000110011001",  "000000000110001101",  "000000000110000000",  "000000000101110100",  "000000000101101000",  "000000000101011100",  "000000000101001111",  "000000000101000011",  "000000000100110111",  "000000000100101010",  "000000000100011110",  "000000000100010010",  "000000000100000101",  "000000000011111001",  "000000000011101100",  "000000000011100000",  "000000000011010100",  "000000000011000111",  "000000000010111011",  "000000000010101110",  "000000000010100010",  "000000000010010110",  "000000000010001001",  "000000000001111101",  "000000000001110000",  "000000000001100100",  "000000000001010111",  "000000000001001011",  "000000000000111110",  "000000000000110010",  "000000000000100101",  "000000000000011001",  "000000000000001100"),("000000000000000000",  "111111111111110100",  "111111111111100111",  "111111111111011011",  "111111111111001110",  "111111111111000001",  "111111111110110101",  "111111111110101000",  "111111111110011100",  "111111111110001111",  "111111111110000011",  "111111111101110110",  "111111111101101010",  "111111111101011101",  "111111111101010001",  "111111111101000100",  "111111111100111000",  "111111111100101011",  "111111111100011111",  "111111111100010010",  "111111111100000101",  "111111111011111001",  "111111111011101100",  "111111111011100000",  "111111111011010011",  "111111111011000111",  "111111111010111010",  "111111111010101101",  "111111111010100001",  "111111111010010100",  "111111111010001000",  "111111111001111011",  "111111111001101111",  "111111111001100010",  "111111111001010101",  "111111111001001001",  "111111111000111100",  "111111111000110000",  "111111111000100011",  "111111111000010110",  "111111111000001010",  "111111110111111101",  "111111110111110001",  "111111110111100100",  "111111110111011000",  "111111110111001011",  "111111110110111110",  "111111110110110010",  "111111110110100101",  "111111110110011001",  "111111110110001100",  "111111110110000000",  "111111110101110011",  "111111110101100110",  "111111110101011010",  "111111110101001101",  "111111110101000001",  "111111110100110100",  "111111110100101000",  "111111110100011011",  "111111110100001110",  "111111110100000010",  "111111110011110101",  "111111110011101001",  "111111110011011100",  "111111110011010000",  "111111110011000011",  "111111110010110111",  "111111110010101010",  "111111110010011110",  "111111110010010001",  "111111110010000101",  "111111110001111000",  "111111110001101011",  "111111110001011111",  "111111110001010010",  "111111110001000110",  "111111110000111001",  "111111110000101101",  "111111110000100000",  "111111110000010100",  "111111110000001000",  "111111101111111011",  "111111101111101111",  "111111101111100010",  "111111101111010110",  "111111101111001001",  "111111101110111101",  "111111101110110000",  "111111101110100100",  "111111101110010111",  "111111101110001011",  "111111101101111111",  "111111101101110010",  "111111101101100110",  "111111101101011001",  "111111101101001101",  "111111101101000001",  "111111101100110100",  "111111101100101000",  "111111101100011011",  "111111101100001111",  "111111101100000011",  "111111101011110110",  "111111101011101010",  "111111101011011110",  "111111101011010001",  "111111101011000101",  "111111101010111001",  "111111101010101101",  "111111101010100000",  "111111101010010100",  "111111101010001000",  "111111101001111011",  "111111101001101111",  "111111101001100011",  "111111101001010111",  "111111101001001010",  "111111101000111110",  "111111101000110010",  "111111101000100110",  "111111101000011010",  "111111101000001110",  "111111101000000001",  "111111100111110101",  "111111100111101001",  "111111100111011101",  "111111100111010001",  "111111100111000101",  "111111100110111001",  "111111100110101100",  "111111100110100000",  "111111100110010100",  "111111100110001000",  "111111100101111100",  "111111100101110000",  "111111100101100100",  "111111100101011000",  "111111100101001100",  "111111100101000000",  "111111100100110100",  "111111100100101000",  "111111100100011100",  "111111100100010000",  "111111100100000100",  "111111100011111000",  "111111100011101100",  "111111100011100001",  "111111100011010101",  "111111100011001001",  "111111100010111101",  "111111100010110001",  "111111100010100101",  "111111100010011010",  "111111100010001110",  "111111100010000010",  "111111100001110110",  "111111100001101010",  "111111100001011111",  "111111100001010011",  "111111100001000111",  "111111100000111011",  "111111100000110000",  "111111100000100100",  "111111100000011000",  "111111100000001101",  "111111100000000001",  "111111011111110110",  "111111011111101010",  "111111011111011110",  "111111011111010011",  "111111011111000111",  "111111011110111100",  "111111011110110000",  "111111011110100101",  "111111011110011001",  "111111011110001110",  "111111011110000010",  "111111011101110111",  "111111011101101011",  "111111011101100000",  "111111011101010101",  "111111011101001001",  "111111011100111110",  "111111011100110010",  "111111011100100111",  "111111011100011100",  "111111011100010001",  "111111011100000101",  "111111011011111010",  "111111011011101111",  "111111011011100100",  "111111011011011000",  "111111011011001101",  "111111011011000010",  "111111011010110111",  "111111011010101100",  "111111011010100001",  "111111011010010110",  "111111011010001010",  "111111011001111111",  "111111011001110100",  "111111011001101001",  "111111011001011110",  "111111011001010011",  "111111011001001000",  "111111011000111101",  "111111011000110011",  "111111011000101000",  "111111011000011101",  "111111011000010010",  "111111011000000111",  "111111010111111100",  "111111010111110001",  "111111010111100111",  "111111010111011100",  "111111010111010001",  "111111010111000110",  "111111010110111100",  "111111010110110001",  "111111010110100110",  "111111010110011100",  "111111010110010001",  "111111010110000111",  "111111010101111100",  "111111010101110001",  "111111010101100111",  "111111010101011100",  "111111010101010010",  "111111010101000111",  "111111010100111101",  "111111010100110011",  "111111010100101000",  "111111010100011110",  "111111010100010011",  "111111010100001001",  "111111010011111111",  "111111010011110100",  "111111010011101010",  "111111010011100000",  "111111010011010110",  "111111010011001100",  "111111010011000001",  "111111010010110111",  "111111010010101101",  "111111010010100011",  "111111010010011001",  "111111010010001111",  "111111010010000101",  "111111010001111011",  "111111010001110001",  "111111010001100111",  "111111010001011101",  "111111010001010011",  "111111010001001001",  "111111010000111111",  "111111010000110110",  "111111010000101100",  "111111010000100010",  "111111010000011000",  "111111010000001110",  "111111010000000101",  "111111001111111011",  "111111001111110001",  "111111001111101000",  "111111001111011110",  "111111001111010101",  "111111001111001011",  "111111001111000001",  "111111001110111000",  "111111001110101111",  "111111001110100101",  "111111001110011100",  "111111001110010010",  "111111001110001001",  "111111001110000000",  "111111001101110110",  "111111001101101101",  "111111001101100100",  "111111001101011010",  "111111001101010001",  "111111001101001000",  "111111001100111111",  "111111001100110110",  "111111001100101101",  "111111001100100100",  "111111001100011011",  "111111001100010010",  "111111001100001001",  "111111001100000000",  "111111001011110111",  "111111001011101110",  "111111001011100101",  "111111001011011100",  "111111001011010011",  "111111001011001010",  "111111001011000010",  "111111001010111001",  "111111001010110000",  "111111001010101000",  "111111001010011111",  "111111001010010110",  "111111001010001110",  "111111001010000101",  "111111001001111101",  "111111001001110100",  "111111001001101100",  "111111001001100011",  "111111001001011011",  "111111001001010010",  "111111001001001010",  "111111001001000010",  "111111001000111001",  "111111001000110001",  "111111001000101001",  "111111001000100001",  "111111001000011001",  "111111001000010000",  "111111001000001000",  "111111001000000000",  "111111000111111000",  "111111000111110000",  "111111000111101000",  "111111000111100000",  "111111000111011000",  "111111000111010000",  "111111000111001001",  "111111000111000001",  "111111000110111001",  "111111000110110001",  "111111000110101001",  "111111000110100010",  "111111000110011010",  "111111000110010010",  "111111000110001011",  "111111000110000011",  "111111000101111100",  "111111000101110100",  "111111000101101101",  "111111000101100101",  "111111000101011110",  "111111000101010110",  "111111000101001111",  "111111000101001000",  "111111000101000001",  "111111000100111001",  "111111000100110010",  "111111000100101011",  "111111000100100100",  "111111000100011101",  "111111000100010110",  "111111000100001110",  "111111000100000111",  "111111000100000000",  "111111000011111010",  "111111000011110011",  "111111000011101100",  "111111000011100101",  "111111000011011110",  "111111000011010111",  "111111000011010001",  "111111000011001010",  "111111000011000011",  "111111000010111101",  "111111000010110110",  "111111000010101111",  "111111000010101001",  "111111000010100010",  "111111000010011100",  "111111000010010101",  "111111000010001111",  "111111000010001001",  "111111000010000010",  "111111000001111100",  "111111000001110110",  "111111000001110000",  "111111000001101001",  "111111000001100011",  "111111000001011101",  "111111000001010111",  "111111000001010001",  "111111000001001011",  "111111000001000101",  "111111000000111111",  "111111000000111001",  "111111000000110011",  "111111000000101101",  "111111000000101000",  "111111000000100010",  "111111000000011100",  "111111000000010110",  "111111000000010001",  "111111000000001011",  "111111000000000110",  "111111000000000000",  "111110111111111011",  "111110111111110101",  "111110111111110000",  "111110111111101010",  "111110111111100101",  "111110111111100000",  "111110111111011010",  "111110111111010101",  "111110111111010000",  "111110111111001011",  "111110111111000101",  "111110111111000000",  "111110111110111011",  "111110111110110110",  "111110111110110001",  "111110111110101100",  "111110111110100111",  "111110111110100011",  "111110111110011110",  "111110111110011001",  "111110111110010100",  "111110111110001111",  "111110111110001011",  "111110111110000110",  "111110111110000010",  "111110111101111101",  "111110111101111000",  "111110111101110100",  "111110111101101111",  "111110111101101011",  "111110111101100111",  "111110111101100010",  "111110111101011110",  "111110111101011010",  "111110111101010110",  "111110111101010001",  "111110111101001101",  "111110111101001001",  "111110111101000101",  "111110111101000001",  "111110111100111101",  "111110111100111001",  "111110111100110101",  "111110111100110001",  "111110111100101101",  "111110111100101010",  "111110111100100110",  "111110111100100010",  "111110111100011111",  "111110111100011011",  "111110111100010111",  "111110111100010100",  "111110111100010000",  "111110111100001101",  "111110111100001001",  "111110111100000110",  "111110111100000011",  "111110111011111111",  "111110111011111100",  "111110111011111001",  "111110111011110101",  "111110111011110010",  "111110111011101111",  "111110111011101100",  "111110111011101001",  "111110111011100110",  "111110111011100011",  "111110111011100000",  "111110111011011101",  "111110111011011010",  "111110111011011000",  "111110111011010101",  "111110111011010010",  "111110111011010000",  "111110111011001101",  "111110111011001010",  "111110111011001000",  "111110111011000101",  "111110111011000011",  "111110111011000000",  "111110111010111110",  "111110111010111100",  "111110111010111001",  "111110111010110111",  "111110111010110101",  "111110111010110011",  "111110111010110000",  "111110111010101110",  "111110111010101100",  "111110111010101010",  "111110111010101000",  "111110111010100110",  "111110111010100100",  "111110111010100011",  "111110111010100001",  "111110111010011111",  "111110111010011101",  "111110111010011011",  "111110111010011010",  "111110111010011000",  "111110111010010111",  "111110111010010101",  "111110111010010100",  "111110111010010010",  "111110111010010001",  "111110111010001111",  "111110111010001110",  "111110111010001101",  "111110111010001100",  "111110111010001010",  "111110111010001001",  "111110111010001000",  "111110111010000111",  "111110111010000110",  "111110111010000101",  "111110111010000100",  "111110111010000011",  "111110111010000010",  "111110111010000001",  "111110111010000001",  "111110111010000000",  "111110111001111111",  "111110111001111111",  "111110111001111110",  "111110111001111101",  "111110111001111101",  "111110111001111100",  "111110111001111100",  "111110111001111100",  "111110111001111011",  "111110111001111011",  "111110111001111011",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111011",  "111110111001111011",  "111110111001111011",  "111110111001111100",  "111110111001111100",  "111110111001111101",  "111110111001111101",  "111110111001111110",  "111110111001111110",  "111110111001111111",  "111110111001111111",  "111110111010000000",  "111110111010000001",  "111110111010000010",  "111110111010000010",  "111110111010000011",  "111110111010000100",  "111110111010000101",  "111110111010000110",  "111110111010000111",  "111110111010001000",  "111110111010001001",  "111110111010001011",  "111110111010001100",  "111110111010001101",  "111110111010001110",  "111110111010010000",  "111110111010010001",  "111110111010010011",  "111110111010010100",  "111110111010010110",  "111110111010010111",  "111110111010011001",  "111110111010011010",  "111110111010011100",  "111110111010011110",  "111110111010100000",  "111110111010100001",  "111110111010100011",  "111110111010100101",  "111110111010100111",  "111110111010101001",  "111110111010101011",  "111110111010101101",  "111110111010101111",  "111110111010110001",  "111110111010110100",  "111110111010110110",  "111110111010111000",  "111110111010111010",  "111110111010111101",  "111110111010111111",  "111110111011000010",  "111110111011000100",  "111110111011000111",  "111110111011001001",  "111110111011001100",  "111110111011001111",  "111110111011010001",  "111110111011010100",  "111110111011010111",  "111110111011011010",  "111110111011011100",  "111110111011011111",  "111110111011100010",  "111110111011100101",  "111110111011101000",  "111110111011101011",  "111110111011101111",  "111110111011110010",  "111110111011110101",  "111110111011111000",  "111110111011111100",  "111110111011111111",  "111110111100000010",  "111110111100000110",  "111110111100001001",  "111110111100001101",  "111110111100010000",  "111110111100010100",  "111110111100010111",  "111110111100011011",  "111110111100011111",  "111110111100100011",  "111110111100100110",  "111110111100101010",  "111110111100101110",  "111110111100110010",  "111110111100110110",  "111110111100111010",  "111110111100111110",  "111110111101000010",  "111110111101000110",  "111110111101001011",  "111110111101001111",  "111110111101010011",  "111110111101010111",  "111110111101011100",  "111110111101100000",  "111110111101100101",  "111110111101101001",  "111110111101101110",  "111110111101110010",  "111110111101110111",  "111110111101111011",  "111110111110000000",  "111110111110000101",  "111110111110001010",  "111110111110001110",  "111110111110010011",  "111110111110011000",  "111110111110011101",  "111110111110100010",  "111110111110100111",  "111110111110101100",  "111110111110110001",  "111110111110110110",  "111110111110111100",  "111110111111000001",  "111110111111000110",  "111110111111001011",  "111110111111010001",  "111110111111010110",  "111110111111011100",  "111110111111100001",  "111110111111100111",  "111110111111101100",  "111110111111110010",  "111110111111110111",  "111110111111111101",  "111111000000000011",  "111111000000001001",  "111111000000001110",  "111111000000010100",  "111111000000011010",  "111111000000100000",  "111111000000100110",  "111111000000101100",  "111111000000110010",  "111111000000111000",  "111111000000111110",  "111111000001000100",  "111111000001001011",  "111111000001010001",  "111111000001010111",  "111111000001011110",  "111111000001100100",  "111111000001101010",  "111111000001110001",  "111111000001110111",  "111111000001111110",  "111111000010000100",  "111111000010001011",  "111111000010010010",  "111111000010011000",  "111111000010011111",  "111111000010100110",  "111111000010101101",  "111111000010110011",  "111111000010111010",  "111111000011000001",  "111111000011001000",  "111111000011001111",  "111111000011010110",  "111111000011011101",  "111111000011100100",  "111111000011101100",  "111111000011110011",  "111111000011111010",  "111111000100000001",  "111111000100001001",  "111111000100010000",  "111111000100010111",  "111111000100011111",  "111111000100100110",  "111111000100101110",  "111111000100110101",  "111111000100111101",  "111111000101000101",  "111111000101001100",  "111111000101010100",  "111111000101011100",  "111111000101100100",  "111111000101101011",  "111111000101110011",  "111111000101111011",  "111111000110000011",  "111111000110001011",  "111111000110010011",  "111111000110011011",  "111111000110100011",  "111111000110101011",  "111111000110110011",  "111111000110111100",  "111111000111000100",  "111111000111001100",  "111111000111010100",  "111111000111011101",  "111111000111100101",  "111111000111101110",  "111111000111110110",  "111111000111111111",  "111111001000000111",  "111111001000010000",  "111111001000011000",  "111111001000100001",  "111111001000101010",  "111111001000110010",  "111111001000111011",  "111111001001000100",  "111111001001001101",  "111111001001010110",  "111111001001011110",  "111111001001100111",  "111111001001110000",  "111111001001111001",  "111111001010000010",  "111111001010001100",  "111111001010010101",  "111111001010011110",  "111111001010100111",  "111111001010110000",  "111111001010111010",  "111111001011000011",  "111111001011001100",  "111111001011010110",  "111111001011011111",  "111111001011101000",  "111111001011110010",  "111111001011111011",  "111111001100000101",  "111111001100001110",  "111111001100011000",  "111111001100100010",  "111111001100101011",  "111111001100110101",  "111111001100111111",  "111111001101001001",  "111111001101010011",  "111111001101011100",  "111111001101100110",  "111111001101110000",  "111111001101111010",  "111111001110000100",  "111111001110001110",  "111111001110011000",  "111111001110100010",  "111111001110101100",  "111111001110110111",  "111111001111000001",  "111111001111001011",  "111111001111010101",  "111111001111100000",  "111111001111101010",  "111111001111110100",  "111111001111111111",  "111111010000001001",  "111111010000010100",  "111111010000011110",  "111111010000101001",  "111111010000110011",  "111111010000111110",  "111111010001001000",  "111111010001010011",  "111111010001011110",  "111111010001101000",  "111111010001110011",  "111111010001111110",  "111111010010001001",  "111111010010010100",  "111111010010011111",  "111111010010101001",  "111111010010110100",  "111111010010111111",  "111111010011001010",  "111111010011010101",  "111111010011100001",  "111111010011101100",  "111111010011110111",  "111111010100000010",  "111111010100001101",  "111111010100011000",  "111111010100100100",  "111111010100101111",  "111111010100111010",  "111111010101000110",  "111111010101010001",  "111111010101011100",  "111111010101101000",  "111111010101110011",  "111111010101111111",  "111111010110001010",  "111111010110010110",  "111111010110100001",  "111111010110101101",  "111111010110111001",  "111111010111000100",  "111111010111010000",  "111111010111011100",  "111111010111101000",  "111111010111110011",  "111111010111111111",  "111111011000001011",  "111111011000010111",  "111111011000100011",  "111111011000101111",  "111111011000111011",  "111111011001000111",  "111111011001010011",  "111111011001011111",  "111111011001101011",  "111111011001110111",  "111111011010000011",  "111111011010001111",  "111111011010011011",  "111111011010101000",  "111111011010110100",  "111111011011000000",  "111111011011001100",  "111111011011011001",  "111111011011100101",  "111111011011110001",  "111111011011111110",  "111111011100001010",  "111111011100010111",  "111111011100100011",  "111111011100110000",  "111111011100111100",  "111111011101001001",  "111111011101010101",  "111111011101100010",  "111111011101101111",  "111111011101111011",  "111111011110001000",  "111111011110010101",  "111111011110100001",  "111111011110101110",  "111111011110111011",  "111111011111001000",  "111111011111010101",  "111111011111100001",  "111111011111101110",  "111111011111111011",  "111111100000001000",  "111111100000010101",  "111111100000100010",  "111111100000101111",  "111111100000111100",  "111111100001001001",  "111111100001010110",  "111111100001100011",  "111111100001110001",  "111111100001111110",  "111111100010001011",  "111111100010011000",  "111111100010100101",  "111111100010110011",  "111111100011000000",  "111111100011001101",  "111111100011011010",  "111111100011101000",  "111111100011110101",  "111111100100000010",  "111111100100010000",  "111111100100011101",  "111111100100101011",  "111111100100111000",  "111111100101000110",  "111111100101010011",  "111111100101100001",  "111111100101101110",  "111111100101111100",  "111111100110001001",  "111111100110010111",  "111111100110100101",  "111111100110110010",  "111111100111000000",  "111111100111001110",  "111111100111011011",  "111111100111101001",  "111111100111110111",  "111111101000000101",  "111111101000010010",  "111111101000100000",  "111111101000101110",  "111111101000111100",  "111111101001001010",  "111111101001011000",  "111111101001100110",  "111111101001110011",  "111111101010000001",  "111111101010001111",  "111111101010011101",  "111111101010101011",  "111111101010111001",  "111111101011000111",  "111111101011010110",  "111111101011100100",  "111111101011110010",  "111111101100000000",  "111111101100001110",  "111111101100011100",  "111111101100101010",  "111111101100111000",  "111111101101000111",  "111111101101010101",  "111111101101100011",  "111111101101110001",  "111111101110000000",  "111111101110001110",  "111111101110011100",  "111111101110101010",  "111111101110111001",  "111111101111000111",  "111111101111010101",  "111111101111100100",  "111111101111110010",  "111111110000000001",  "111111110000001111",  "111111110000011101",  "111111110000101100",  "111111110000111010",  "111111110001001001",  "111111110001010111",  "111111110001100110",  "111111110001110100",  "111111110010000011",  "111111110010010001",  "111111110010100000",  "111111110010101111",  "111111110010111101",  "111111110011001100",  "111111110011011010",  "111111110011101001",  "111111110011111000",  "111111110100000110",  "111111110100010101",  "111111110100100100",  "111111110100110010",  "111111110101000001",  "111111110101010000",  "111111110101011111",  "111111110101101101",  "111111110101111100",  "111111110110001011",  "111111110110011010",  "111111110110101000",  "111111110110110111",  "111111110111000110",  "111111110111010101",  "111111110111100100",  "111111110111110011",  "111111111000000001",  "111111111000010000",  "111111111000011111",  "111111111000101110",  "111111111000111101",  "111111111001001100",  "111111111001011011",  "111111111001101010",  "111111111001111001",  "111111111010001000",  "111111111010010111",  "111111111010100110",  "111111111010110101",  "111111111011000100",  "111111111011010010",  "111111111011100010",  "111111111011110001",  "111111111100000000",  "111111111100001111",  "111111111100011110",  "111111111100101101",  "111111111100111100",  "111111111101001011",  "111111111101011010",  "111111111101101001",  "111111111101111000",  "111111111110000111",  "111111111110010110",  "111111111110100101",  "111111111110110100",  "111111111111000011",  "111111111111010011",  "111111111111100010",  "111111111111110001"),("000000000000000000",  "000000000000001111",  "000000000000011110",  "000000000000101101",  "000000000000111101",  "000000000001001100",  "000000000001011011",  "000000000001101010",  "000000000001111001",  "000000000010001001",  "000000000010011000",  "000000000010100111",  "000000000010110110",  "000000000011000101",  "000000000011010101",  "000000000011100100",  "000000000011110011",  "000000000100000010",  "000000000100010001",  "000000000100100001",  "000000000100110000",  "000000000100111111",  "000000000101001110",  "000000000101011110",  "000000000101101101",  "000000000101111100",  "000000000110001011",  "000000000110011011",  "000000000110101010",  "000000000110111001",  "000000000111001000",  "000000000111011000",  "000000000111100111",  "000000000111110110",  "000000001000000101",  "000000001000010101",  "000000001000100100",  "000000001000110011",  "000000001001000010",  "000000001001010010",  "000000001001100001",  "000000001001110000",  "000000001001111111",  "000000001010001111",  "000000001010011110",  "000000001010101101",  "000000001010111100",  "000000001011001100",  "000000001011011011",  "000000001011101010",  "000000001011111001",  "000000001100001001",  "000000001100011000",  "000000001100100111",  "000000001100110111",  "000000001101000110",  "000000001101010101",  "000000001101100100",  "000000001101110100",  "000000001110000011",  "000000001110010010",  "000000001110100001",  "000000001110110000",  "000000001111000000",  "000000001111001111",  "000000001111011110",  "000000001111101101",  "000000001111111101",  "000000010000001100",  "000000010000011011",  "000000010000101010",  "000000010000111001",  "000000010001001001",  "000000010001011000",  "000000010001100111",  "000000010001110110",  "000000010010000101",  "000000010010010101",  "000000010010100100",  "000000010010110011",  "000000010011000010",  "000000010011010001",  "000000010011100000",  "000000010011101111",  "000000010011111111",  "000000010100001110",  "000000010100011101",  "000000010100101100",  "000000010100111011",  "000000010101001010",  "000000010101011001",  "000000010101101000",  "000000010101110111",  "000000010110000110",  "000000010110010110",  "000000010110100101",  "000000010110110100",  "000000010111000011",  "000000010111010010",  "000000010111100001",  "000000010111110000",  "000000010111111111",  "000000011000001110",  "000000011000011101",  "000000011000101100",  "000000011000111011",  "000000011001001010",  "000000011001011001",  "000000011001101000",  "000000011001110111",  "000000011010000101",  "000000011010010100",  "000000011010100011",  "000000011010110010",  "000000011011000001",  "000000011011010000",  "000000011011011111",  "000000011011101110",  "000000011011111100",  "000000011100001011",  "000000011100011010",  "000000011100101001",  "000000011100111000",  "000000011101000111",  "000000011101010101",  "000000011101100100",  "000000011101110011",  "000000011110000010",  "000000011110010000",  "000000011110011111",  "000000011110101110",  "000000011110111100",  "000000011111001011",  "000000011111011010",  "000000011111101000",  "000000011111110111",  "000000100000000110",  "000000100000010100",  "000000100000100011",  "000000100000110001",  "000000100001000000",  "000000100001001110",  "000000100001011101",  "000000100001101100",  "000000100001111010",  "000000100010001001",  "000000100010010111",  "000000100010100101",  "000000100010110100",  "000000100011000010",  "000000100011010001",  "000000100011011111",  "000000100011101110",  "000000100011111100",  "000000100100001010",  "000000100100011001",  "000000100100100111",  "000000100100110101",  "000000100101000100",  "000000100101010010",  "000000100101100000",  "000000100101101110",  "000000100101111100",  "000000100110001011",  "000000100110011001",  "000000100110100111",  "000000100110110101",  "000000100111000011",  "000000100111010001",  "000000100111100000",  "000000100111101110",  "000000100111111100",  "000000101000001010",  "000000101000011000",  "000000101000100110",  "000000101000110100",  "000000101001000010",  "000000101001010000",  "000000101001011110",  "000000101001101011",  "000000101001111001",  "000000101010000111",  "000000101010010101",  "000000101010100011",  "000000101010110001",  "000000101010111110",  "000000101011001100",  "000000101011011010",  "000000101011101000",  "000000101011110101",  "000000101100000011",  "000000101100010001",  "000000101100011110",  "000000101100101100",  "000000101100111010",  "000000101101000111",  "000000101101010101",  "000000101101100010",  "000000101101110000",  "000000101101111101",  "000000101110001011",  "000000101110011000",  "000000101110100101",  "000000101110110011",  "000000101111000000",  "000000101111001110",  "000000101111011011",  "000000101111101000",  "000000101111110101",  "000000110000000011",  "000000110000010000",  "000000110000011101",  "000000110000101010",  "000000110000110111",  "000000110001000101",  "000000110001010010",  "000000110001011111",  "000000110001101100",  "000000110001111001",  "000000110010000110",  "000000110010010011",  "000000110010100000",  "000000110010101101",  "000000110010111010",  "000000110011000111",  "000000110011010011",  "000000110011100000",  "000000110011101101",  "000000110011111010",  "000000110100000111",  "000000110100010011",  "000000110100100000",  "000000110100101101",  "000000110100111001",  "000000110101000110",  "000000110101010010",  "000000110101011111",  "000000110101101100",  "000000110101111000",  "000000110110000101",  "000000110110010001",  "000000110110011101",  "000000110110101010",  "000000110110110110",  "000000110111000011",  "000000110111001111",  "000000110111011011",  "000000110111100111",  "000000110111110100",  "000000111000000000",  "000000111000001100",  "000000111000011000",  "000000111000100100",  "000000111000110000",  "000000111000111100",  "000000111001001000",  "000000111001010100",  "000000111001100000",  "000000111001101100",  "000000111001111000",  "000000111010000100",  "000000111010010000",  "000000111010011100",  "000000111010100111",  "000000111010110011",  "000000111010111111",  "000000111011001011",  "000000111011010110",  "000000111011100010",  "000000111011101101",  "000000111011111001",  "000000111100000101",  "000000111100010000",  "000000111100011011",  "000000111100100111",  "000000111100110010",  "000000111100111110",  "000000111101001001",  "000000111101010100",  "000000111101100000",  "000000111101101011",  "000000111101110110",  "000000111110000001",  "000000111110001100",  "000000111110010111",  "000000111110100010",  "000000111110101110",  "000000111110111001",  "000000111111000100",  "000000111111001110",  "000000111111011001",  "000000111111100100",  "000000111111101111",  "000000111111111010",  "000001000000000101",  "000001000000001111",  "000001000000011010",  "000001000000100101",  "000001000000101111",  "000001000000111010",  "000001000001000100",  "000001000001001111",  "000001000001011001",  "000001000001100100",  "000001000001101110",  "000001000001111001",  "000001000010000011",  "000001000010001101",  "000001000010011000",  "000001000010100010",  "000001000010101100",  "000001000010110110",  "000001000011000000",  "000001000011001010",  "000001000011010101",  "000001000011011111",  "000001000011101001",  "000001000011110010",  "000001000011111100",  "000001000100000110",  "000001000100010000",  "000001000100011010",  "000001000100100100",  "000001000100101101",  "000001000100110111",  "000001000101000001",  "000001000101001010",  "000001000101010100",  "000001000101011101",  "000001000101100111",  "000001000101110000",  "000001000101111010",  "000001000110000011",  "000001000110001101",  "000001000110010110",  "000001000110011111",  "000001000110101000",  "000001000110110001",  "000001000110111011",  "000001000111000100",  "000001000111001101",  "000001000111010110",  "000001000111011111",  "000001000111101000",  "000001000111110001",  "000001000111111010",  "000001001000000010",  "000001001000001011",  "000001001000010100",  "000001001000011101",  "000001001000100101",  "000001001000101110",  "000001001000110110",  "000001001000111111",  "000001001001001000",  "000001001001010000",  "000001001001011000",  "000001001001100001",  "000001001001101001",  "000001001001110001",  "000001001001111010",  "000001001010000010",  "000001001010001010",  "000001001010010010",  "000001001010011010",  "000001001010100010",  "000001001010101010",  "000001001010110010",  "000001001010111010",  "000001001011000010",  "000001001011001010",  "000001001011010010",  "000001001011011010",  "000001001011100001",  "000001001011101001",  "000001001011110001",  "000001001011111000",  "000001001100000000",  "000001001100000111",  "000001001100001111",  "000001001100010110",  "000001001100011101",  "000001001100100101",  "000001001100101100",  "000001001100110011",  "000001001100111010",  "000001001101000010",  "000001001101001001",  "000001001101010000",  "000001001101010111",  "000001001101011110",  "000001001101100101",  "000001001101101100",  "000001001101110010",  "000001001101111001",  "000001001110000000",  "000001001110000111",  "000001001110001101",  "000001001110010100",  "000001001110011011",  "000001001110100001",  "000001001110101000",  "000001001110101110",  "000001001110110100",  "000001001110111011",  "000001001111000001",  "000001001111000111",  "000001001111001110",  "000001001111010100",  "000001001111011010",  "000001001111100000",  "000001001111100110",  "000001001111101100",  "000001001111110010",  "000001001111111000",  "000001001111111110",  "000001010000000100",  "000001010000001001",  "000001010000001111",  "000001010000010101",  "000001010000011010",  "000001010000100000",  "000001010000100101",  "000001010000101011",  "000001010000110000",  "000001010000110110",  "000001010000111011",  "000001010001000000",  "000001010001000110",  "000001010001001011",  "000001010001010000",  "000001010001010101",  "000001010001011010",  "000001010001011111",  "000001010001100100",  "000001010001101001",  "000001010001101110",  "000001010001110011",  "000001010001111000",  "000001010001111100",  "000001010010000001",  "000001010010000110",  "000001010010001010",  "000001010010001111",  "000001010010010011",  "000001010010011000",  "000001010010011100",  "000001010010100000",  "000001010010100101",  "000001010010101001",  "000001010010101101",  "000001010010110001",  "000001010010110101",  "000001010010111001",  "000001010010111101",  "000001010011000001",  "000001010011000101",  "000001010011001001",  "000001010011001101",  "000001010011010001",  "000001010011010101",  "000001010011011000",  "000001010011011100",  "000001010011011111",  "000001010011100011",  "000001010011100110",  "000001010011101010",  "000001010011101101",  "000001010011110000",  "000001010011110100",  "000001010011110111",  "000001010011111010",  "000001010011111101",  "000001010100000000",  "000001010100000011",  "000001010100000110",  "000001010100001001",  "000001010100001100",  "000001010100001111",  "000001010100010010",  "000001010100010101",  "000001010100010111",  "000001010100011010",  "000001010100011100",  "000001010100011111",  "000001010100100001",  "000001010100100100",  "000001010100100110",  "000001010100101001",  "000001010100101011",  "000001010100101101",  "000001010100101111",  "000001010100110001",  "000001010100110011",  "000001010100110110",  "000001010100110111",  "000001010100111001",  "000001010100111011",  "000001010100111101",  "000001010100111111",  "000001010101000001",  "000001010101000010",  "000001010101000100",  "000001010101000101",  "000001010101000111",  "000001010101001000",  "000001010101001010",  "000001010101001011",  "000001010101001101",  "000001010101001110",  "000001010101001111",  "000001010101010000",  "000001010101010001",  "000001010101010010",  "000001010101010011",  "000001010101010100",  "000001010101010101",  "000001010101010110",  "000001010101010111",  "000001010101011000",  "000001010101011000",  "000001010101011001",  "000001010101011010",  "000001010101011010",  "000001010101011011",  "000001010101011011",  "000001010101011100",  "000001010101011100",  "000001010101011100",  "000001010101011100",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011100",  "000001010101011100",  "000001010101011100",  "000001010101011011",  "000001010101011011",  "000001010101011010",  "000001010101011010",  "000001010101011001",  "000001010101011001",  "000001010101011000",  "000001010101010111",  "000001010101010111",  "000001010101010110",  "000001010101010101",  "000001010101010100",  "000001010101010011",  "000001010101010010",  "000001010101010001",  "000001010101010000",  "000001010101001110",  "000001010101001101",  "000001010101001100",  "000001010101001010",  "000001010101001001",  "000001010101001000",  "000001010101000110",  "000001010101000100",  "000001010101000011",  "000001010101000001",  "000001010100111111",  "000001010100111110",  "000001010100111100",  "000001010100111010",  "000001010100111000",  "000001010100110110",  "000001010100110100",  "000001010100110010",  "000001010100110000",  "000001010100101110",  "000001010100101011",  "000001010100101001",  "000001010100100111",  "000001010100100100",  "000001010100100010",  "000001010100011111",  "000001010100011101",  "000001010100011010",  "000001010100010111",  "000001010100010101",  "000001010100010010",  "000001010100001111",  "000001010100001100",  "000001010100001001",  "000001010100000110",  "000001010100000011",  "000001010100000000",  "000001010011111101",  "000001010011111010",  "000001010011110111",  "000001010011110011",  "000001010011110000",  "000001010011101101",  "000001010011101001",  "000001010011100110",  "000001010011100010",  "000001010011011111",  "000001010011011011",  "000001010011010111",  "000001010011010011",  "000001010011010000",  "000001010011001100",  "000001010011001000",  "000001010011000100",  "000001010011000000",  "000001010010111100",  "000001010010111000",  "000001010010110100",  "000001010010101111",  "000001010010101011",  "000001010010100111",  "000001010010100010",  "000001010010011110",  "000001010010011001",  "000001010010010101",  "000001010010010000",  "000001010010001100",  "000001010010000111",  "000001010010000010",  "000001010001111110",  "000001010001111001",  "000001010001110100",  "000001010001101111",  "000001010001101010",  "000001010001100101",  "000001010001100000",  "000001010001011011",  "000001010001010101",  "000001010001010000",  "000001010001001011",  "000001010001000101",  "000001010001000000",  "000001010000111011",  "000001010000110101",  "000001010000110000",  "000001010000101010",  "000001010000100100",  "000001010000011111",  "000001010000011001",  "000001010000010011",  "000001010000001101",  "000001010000000111",  "000001010000000001",  "000001001111111011",  "000001001111110101",  "000001001111101111",  "000001001111101001",  "000001001111100011",  "000001001111011100",  "000001001111010110",  "000001001111010000",  "000001001111001001",  "000001001111000011",  "000001001110111100",  "000001001110110110",  "000001001110101111",  "000001001110101000",  "000001001110100010",  "000001001110011011",  "000001001110010100",  "000001001110001101",  "000001001110000110",  "000001001101111111",  "000001001101111000",  "000001001101110001",  "000001001101101010",  "000001001101100011",  "000001001101011100",  "000001001101010101",  "000001001101001101",  "000001001101000110",  "000001001100111110",  "000001001100110111",  "000001001100101111",  "000001001100101000",  "000001001100100000",  "000001001100011001",  "000001001100010001",  "000001001100001001",  "000001001100000001",  "000001001011111001",  "000001001011110010",  "000001001011101010",  "000001001011100010",  "000001001011011001",  "000001001011010001",  "000001001011001001",  "000001001011000001",  "000001001010111001",  "000001001010110000",  "000001001010101000",  "000001001010100000",  "000001001010010111",  "000001001010001111",  "000001001010000110",  "000001001001111110",  "000001001001110101",  "000001001001101100",  "000001001001100100",  "000001001001011011",  "000001001001010010",  "000001001001001001",  "000001001001000000",  "000001001000110111",  "000001001000101110",  "000001001000100101",  "000001001000011100",  "000001001000010011",  "000001001000001010",  "000001001000000000",  "000001000111110111",  "000001000111101110",  "000001000111100100",  "000001000111011011",  "000001000111010001",  "000001000111001000",  "000001000110111110",  "000001000110110101",  "000001000110101011",  "000001000110100001",  "000001000110010111",  "000001000110001110",  "000001000110000100",  "000001000101111010",  "000001000101110000",  "000001000101100110",  "000001000101011100",  "000001000101010010",  "000001000101000111",  "000001000100111101",  "000001000100110011",  "000001000100101001",  "000001000100011110",  "000001000100010100",  "000001000100001010",  "000001000011111111",  "000001000011110101",  "000001000011101010",  "000001000011011111",  "000001000011010101",  "000001000011001010",  "000001000010111111",  "000001000010110101",  "000001000010101010",  "000001000010011111",  "000001000010010100",  "000001000010001001",  "000001000001111110",  "000001000001110011",  "000001000001101000",  "000001000001011101",  "000001000001010010",  "000001000001000110",  "000001000000111011",  "000001000000110000",  "000001000000100100",  "000001000000011001",  "000001000000001110",  "000001000000000010",  "000000111111110111",  "000000111111101011",  "000000111111011111",  "000000111111010100",  "000000111111001000",  "000000111110111100",  "000000111110110000",  "000000111110100101",  "000000111110011001",  "000000111110001101",  "000000111110000001",  "000000111101110101",  "000000111101101001",  "000000111101011101",  "000000111101010001",  "000000111101000100",  "000000111100111000",  "000000111100101100",  "000000111100100000",  "000000111100010011",  "000000111100000111",  "000000111011111011",  "000000111011101110",  "000000111011100010",  "000000111011010101",  "000000111011001000",  "000000111010111100",  "000000111010101111",  "000000111010100010",  "000000111010010110",  "000000111010001001",  "000000111001111100",  "000000111001101111",  "000000111001100010",  "000000111001010101",  "000000111001001000",  "000000111000111011",  "000000111000101110",  "000000111000100001",  "000000111000010100",  "000000111000000111",  "000000110111111010",  "000000110111101100",  "000000110111011111",  "000000110111010010",  "000000110111000100",  "000000110110110111",  "000000110110101001",  "000000110110011100",  "000000110110001110",  "000000110110000001",  "000000110101110011",  "000000110101100110",  "000000110101011000",  "000000110101001010",  "000000110100111100",  "000000110100101111",  "000000110100100001",  "000000110100010011",  "000000110100000101",  "000000110011110111",  "000000110011101001",  "000000110011011011",  "000000110011001101",  "000000110010111111",  "000000110010110001",  "000000110010100011",  "000000110010010100",  "000000110010000110",  "000000110001111000",  "000000110001101010",  "000000110001011011",  "000000110001001101",  "000000110000111110",  "000000110000110000",  "000000110000100001",  "000000110000010011",  "000000110000000100",  "000000101111110110",  "000000101111100111",  "000000101111011000",  "000000101111001010",  "000000101110111011",  "000000101110101100",  "000000101110011101",  "000000101110001111",  "000000101110000000",  "000000101101110001",  "000000101101100010",  "000000101101010011",  "000000101101000100",  "000000101100110101",  "000000101100100110",  "000000101100010111",  "000000101100000111",  "000000101011111000",  "000000101011101001",  "000000101011011010",  "000000101011001011",  "000000101010111011",  "000000101010101100",  "000000101010011101",  "000000101010001101",  "000000101001111110",  "000000101001101110",  "000000101001011111",  "000000101001001111",  "000000101001000000",  "000000101000110000",  "000000101000100000",  "000000101000010001",  "000000101000000001",  "000000100111110001",  "000000100111100010",  "000000100111010010",  "000000100111000010",  "000000100110110010",  "000000100110100010",  "000000100110010011",  "000000100110000011",  "000000100101110011",  "000000100101100011",  "000000100101010011",  "000000100101000011",  "000000100100110011",  "000000100100100010",  "000000100100010010",  "000000100100000010",  "000000100011110010",  "000000100011100010",  "000000100011010001",  "000000100011000001",  "000000100010110001",  "000000100010100001",  "000000100010010000",  "000000100010000000",  "000000100001101111",  "000000100001011111",  "000000100001001111",  "000000100000111110",  "000000100000101110",  "000000100000011101",  "000000100000001100",  "000000011111111100",  "000000011111101011",  "000000011111011011",  "000000011111001010",  "000000011110111001",  "000000011110101000",  "000000011110011000",  "000000011110000111",  "000000011101110110",  "000000011101100101",  "000000011101010100",  "000000011101000100",  "000000011100110011",  "000000011100100010",  "000000011100010001",  "000000011100000000",  "000000011011101111",  "000000011011011110",  "000000011011001101",  "000000011010111100",  "000000011010101011",  "000000011010011010",  "000000011010001000",  "000000011001110111",  "000000011001100110",  "000000011001010101",  "000000011001000100",  "000000011000110010",  "000000011000100001",  "000000011000010000",  "000000010111111111",  "000000010111101101",  "000000010111011100",  "000000010111001010",  "000000010110111001",  "000000010110101000",  "000000010110010110",  "000000010110000101",  "000000010101110011",  "000000010101100010",  "000000010101010000",  "000000010100111111",  "000000010100101101",  "000000010100011100",  "000000010100001010",  "000000010011111000",  "000000010011100111",  "000000010011010101",  "000000010011000011",  "000000010010110010",  "000000010010100000",  "000000010010001110",  "000000010001111100",  "000000010001101011",  "000000010001011001",  "000000010001000111",  "000000010000110101",  "000000010000100011",  "000000010000010010",  "000000010000000000",  "000000001111101110",  "000000001111011100",  "000000001111001010",  "000000001110111000",  "000000001110100110",  "000000001110010100",  "000000001110000010",  "000000001101110000",  "000000001101011110",  "000000001101001100",  "000000001100111010",  "000000001100101000",  "000000001100010110",  "000000001100000100",  "000000001011110001",  "000000001011011111",  "000000001011001101",  "000000001010111011",  "000000001010101001",  "000000001010010111",  "000000001010000100",  "000000001001110010",  "000000001001100000",  "000000001001001110",  "000000001000111100",  "000000001000101001",  "000000001000010111",  "000000001000000101",  "000000000111110010",  "000000000111100000",  "000000000111001110",  "000000000110111011",  "000000000110101001",  "000000000110010111",  "000000000110000100",  "000000000101110010",  "000000000101100000",  "000000000101001101",  "000000000100111011",  "000000000100101000",  "000000000100010110",  "000000000100000011",  "000000000011110001",  "000000000011011110",  "000000000011001100",  "000000000010111001",  "000000000010100111",  "000000000010010100",  "000000000010000010",  "000000000001101111",  "000000000001011101",  "000000000001001010",  "000000000000111000",  "000000000000100101",  "000000000000010011"),("000000000000000000",  "111111111111101101",  "111111111111011011",  "111111111111001000",  "111111111110110110",  "111111111110100011",  "111111111110010000",  "111111111101111110",  "111111111101101011",  "111111111101011000",  "111111111101000110",  "111111111100110011",  "111111111100100000",  "111111111100001110",  "111111111011111011",  "111111111011101000",  "111111111011010110",  "111111111011000011",  "111111111010110000",  "111111111010011110",  "111111111010001011",  "111111111001111000",  "111111111001100110",  "111111111001010011",  "111111111001000000",  "111111111000101101",  "111111111000011011",  "111111111000001000",  "111111110111110101",  "111111110111100011",  "111111110111010000",  "111111110110111101",  "111111110110101010",  "111111110110011000",  "111111110110000101",  "111111110101110010",  "111111110101011111",  "111111110101001101",  "111111110100111010",  "111111110100100111",  "111111110100010100",  "111111110100000010",  "111111110011101111",  "111111110011011100",  "111111110011001001",  "111111110010110110",  "111111110010100100",  "111111110010010001",  "111111110001111110",  "111111110001101011",  "111111110001011001",  "111111110001000110",  "111111110000110011",  "111111110000100000",  "111111110000001110",  "111111101111111011",  "111111101111101000",  "111111101111010101",  "111111101111000011",  "111111101110110000",  "111111101110011101",  "111111101110001011",  "111111101101111000",  "111111101101100101",  "111111101101010010",  "111111101101000000",  "111111101100101101",  "111111101100011010",  "111111101100000111",  "111111101011110101",  "111111101011100010",  "111111101011001111",  "111111101010111101",  "111111101010101010",  "111111101010010111",  "111111101010000101",  "111111101001110010",  "111111101001011111",  "111111101001001101",  "111111101000111010",  "111111101000100111",  "111111101000010101",  "111111101000000010",  "111111100111101111",  "111111100111011101",  "111111100111001010",  "111111100110111000",  "111111100110100101",  "111111100110010010",  "111111100110000000",  "111111100101101101",  "111111100101011011",  "111111100101001000",  "111111100100110110",  "111111100100100011",  "111111100100010000",  "111111100011111110",  "111111100011101011",  "111111100011011001",  "111111100011000110",  "111111100010110100",  "111111100010100001",  "111111100010001111",  "111111100001111101",  "111111100001101010",  "111111100001011000",  "111111100001000101",  "111111100000110011",  "111111100000100000",  "111111100000001110",  "111111011111111100",  "111111011111101001",  "111111011111010111",  "111111011111000101",  "111111011110110010",  "111111011110100000",  "111111011110001110",  "111111011101111011",  "111111011101101001",  "111111011101010111",  "111111011101000100",  "111111011100110010",  "111111011100100000",  "111111011100001110",  "111111011011111100",  "111111011011101001",  "111111011011010111",  "111111011011000101",  "111111011010110011",  "111111011010100001",  "111111011010001111",  "111111011001111101",  "111111011001101010",  "111111011001011000",  "111111011001000110",  "111111011000110100",  "111111011000100010",  "111111011000010000",  "111111010111111110",  "111111010111101100",  "111111010111011010",  "111111010111001000",  "111111010110110110",  "111111010110100101",  "111111010110010011",  "111111010110000001",  "111111010101101111",  "111111010101011101",  "111111010101001011",  "111111010100111010",  "111111010100101000",  "111111010100010110",  "111111010100000100",  "111111010011110011",  "111111010011100001",  "111111010011001111",  "111111010010111101",  "111111010010101100",  "111111010010011010",  "111111010010001001",  "111111010001110111",  "111111010001100101",  "111111010001010100",  "111111010001000010",  "111111010000110001",  "111111010000011111",  "111111010000001110",  "111111001111111101",  "111111001111101011",  "111111001111011010",  "111111001111001000",  "111111001110110111",  "111111001110100110",  "111111001110010100",  "111111001110000011",  "111111001101110010",  "111111001101100001",  "111111001101001111",  "111111001100111110",  "111111001100101101",  "111111001100011100",  "111111001100001011",  "111111001011111010",  "111111001011101001",  "111111001011011000",  "111111001011000111",  "111111001010110110",  "111111001010100101",  "111111001010010100",  "111111001010000011",  "111111001001110010",  "111111001001100001",  "111111001001010000",  "111111001000111111",  "111111001000101110",  "111111001000011110",  "111111001000001101",  "111111000111111100",  "111111000111101100",  "111111000111011011",  "111111000111001010",  "111111000110111010",  "111111000110101001",  "111111000110011001",  "111111000110001000",  "111111000101111000",  "111111000101100111",  "111111000101010111",  "111111000101000110",  "111111000100110110",  "111111000100100101",  "111111000100010101",  "111111000100000101",  "111111000011110101",  "111111000011100100",  "111111000011010100",  "111111000011000100",  "111111000010110100",  "111111000010100100",  "111111000010010100",  "111111000010000100",  "111111000001110100",  "111111000001100100",  "111111000001010100",  "111111000001000100",  "111111000000110100",  "111111000000100100",  "111111000000010100",  "111111000000000100",  "111110111111110101",  "111110111111100101",  "111110111111010101",  "111110111111000101",  "111110111110110110",  "111110111110100110",  "111110111110010111",  "111110111110000111",  "111110111101110111",  "111110111101101000",  "111110111101011001",  "111110111101001001",  "111110111100111010",  "111110111100101010",  "111110111100011011",  "111110111100001100",  "111110111011111101",  "111110111011101101",  "111110111011011110",  "111110111011001111",  "111110111011000000",  "111110111010110001",  "111110111010100010",  "111110111010010011",  "111110111010000100",  "111110111001110101",  "111110111001100110",  "111110111001010111",  "111110111001001000",  "111110111000111010",  "111110111000101011",  "111110111000011100",  "111110111000001110",  "111110110111111111",  "111110110111110000",  "111110110111100010",  "111110110111010011",  "111110110111000101",  "111110110110110110",  "111110110110101000",  "111110110110011010",  "111110110110001011",  "111110110101111101",  "111110110101101111",  "111110110101100000",  "111110110101010010",  "111110110101000100",  "111110110100110110",  "111110110100101000",  "111110110100011010",  "111110110100001100",  "111110110011111110",  "111110110011110000",  "111110110011100010",  "111110110011010100",  "111110110011000111",  "111110110010111001",  "111110110010101011",  "111110110010011110",  "111110110010010000",  "111110110010000010",  "111110110001110101",  "111110110001100111",  "111110110001011010",  "111110110001001101",  "111110110000111111",  "111110110000110010",  "111110110000100101",  "111110110000010111",  "111110110000001010",  "111110101111111101",  "111110101111110000",  "111110101111100011",  "111110101111010110",  "111110101111001001",  "111110101110111100",  "111110101110101111",  "111110101110100010",  "111110101110010101",  "111110101110001001",  "111110101101111100",  "111110101101101111",  "111110101101100011",  "111110101101010110",  "111110101101001001",  "111110101100111101",  "111110101100110000",  "111110101100100100",  "111110101100011000",  "111110101100001011",  "111110101011111111",  "111110101011110011",  "111110101011100111",  "111110101011011011",  "111110101011001110",  "111110101011000010",  "111110101010110110",  "111110101010101010",  "111110101010011111",  "111110101010010011",  "111110101010000111",  "111110101001111011",  "111110101001101111",  "111110101001100100",  "111110101001011000",  "111110101001001101",  "111110101001000001",  "111110101000110110",  "111110101000101010",  "111110101000011111",  "111110101000010011",  "111110101000001000",  "111110100111111101",  "111110100111110010",  "111110100111100110",  "111110100111011011",  "111110100111010000",  "111110100111000101",  "111110100110111010",  "111110100110110000",  "111110100110100101",  "111110100110011010",  "111110100110001111",  "111110100110000100",  "111110100101111010",  "111110100101101111",  "111110100101100101",  "111110100101011010",  "111110100101010000",  "111110100101000101",  "111110100100111011",  "111110100100110001",  "111110100100100110",  "111110100100011100",  "111110100100010010",  "111110100100001000",  "111110100011111110",  "111110100011110100",  "111110100011101010",  "111110100011100000",  "111110100011010110",  "111110100011001100",  "111110100011000011",  "111110100010111001",  "111110100010101111",  "111110100010100110",  "111110100010011100",  "111110100010010011",  "111110100010001001",  "111110100010000000",  "111110100001110111",  "111110100001101101",  "111110100001100100",  "111110100001011011",  "111110100001010010",  "111110100001001001",  "111110100001000000",  "111110100000110111",  "111110100000101110",  "111110100000100101",  "111110100000011100",  "111110100000010100",  "111110100000001011",  "111110100000000010",  "111110011111111010",  "111110011111110001",  "111110011111101001",  "111110011111100000",  "111110011111011000",  "111110011111010000",  "111110011111000111",  "111110011110111111",  "111110011110110111",  "111110011110101111",  "111110011110100111",  "111110011110011111",  "111110011110010111",  "111110011110001111",  "111110011110001000",  "111110011110000000",  "111110011101111000",  "111110011101110000",  "111110011101101001",  "111110011101100001",  "111110011101011010",  "111110011101010010",  "111110011101001011",  "111110011101000100",  "111110011100111101",  "111110011100110101",  "111110011100101110",  "111110011100100111",  "111110011100100000",  "111110011100011001",  "111110011100010010",  "111110011100001100",  "111110011100000101",  "111110011011111110",  "111110011011110111",  "111110011011110001",  "111110011011101010",  "111110011011100100",  "111110011011011101",  "111110011011010111",  "111110011011010001",  "111110011011001010",  "111110011011000100",  "111110011010111110",  "111110011010111000",  "111110011010110010",  "111110011010101100",  "111110011010100110",  "111110011010100000",  "111110011010011010",  "111110011010010101",  "111110011010001111",  "111110011010001001",  "111110011010000100",  "111110011001111110",  "111110011001111001",  "111110011001110011",  "111110011001101110",  "111110011001101001",  "111110011001100100",  "111110011001011110",  "111110011001011001",  "111110011001010100",  "111110011001001111",  "111110011001001010",  "111110011001000110",  "111110011001000001",  "111110011000111100",  "111110011000110111",  "111110011000110011",  "111110011000101110",  "111110011000101010",  "111110011000100101",  "111110011000100001",  "111110011000011101",  "111110011000011001",  "111110011000010100",  "111110011000010000",  "111110011000001100",  "111110011000001000",  "111110011000000100",  "111110011000000000",  "111110010111111101",  "111110010111111001",  "111110010111110101",  "111110010111110001",  "111110010111101110",  "111110010111101010",  "111110010111100111",  "111110010111100100",  "111110010111100000",  "111110010111011101",  "111110010111011010",  "111110010111010111",  "111110010111010100",  "111110010111010001",  "111110010111001110",  "111110010111001011",  "111110010111001000",  "111110010111000101",  "111110010111000010",  "111110010111000000",  "111110010110111101",  "111110010110111011",  "111110010110111000",  "111110010110110110",  "111110010110110100",  "111110010110110001",  "111110010110101111",  "111110010110101101",  "111110010110101011",  "111110010110101001",  "111110010110100111",  "111110010110100101",  "111110010110100011",  "111110010110100001",  "111110010110100000",  "111110010110011110",  "111110010110011101",  "111110010110011011",  "111110010110011010",  "111110010110011000",  "111110010110010111",  "111110010110010110",  "111110010110010100",  "111110010110010011",  "111110010110010010",  "111110010110010001",  "111110010110010000",  "111110010110001111",  "111110010110001111",  "111110010110001110",  "111110010110001101",  "111110010110001100",  "111110010110001100",  "111110010110001011",  "111110010110001011",  "111110010110001011",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001011",  "111110010110001011",  "111110010110001100",  "111110010110001100",  "111110010110001101",  "111110010110001101",  "111110010110001110",  "111110010110001111",  "111110010110010000",  "111110010110010001",  "111110010110010010",  "111110010110010011",  "111110010110010100",  "111110010110010101",  "111110010110010110",  "111110010110010111",  "111110010110011001",  "111110010110011010",  "111110010110011100",  "111110010110011101",  "111110010110011111",  "111110010110100001",  "111110010110100010",  "111110010110100100",  "111110010110100110",  "111110010110101000",  "111110010110101010",  "111110010110101100",  "111110010110101110",  "111110010110110000",  "111110010110110011",  "111110010110110101",  "111110010110110111",  "111110010110111010",  "111110010110111100",  "111110010110111111",  "111110010111000010",  "111110010111000100",  "111110010111000111",  "111110010111001010",  "111110010111001101",  "111110010111010000",  "111110010111010011",  "111110010111010110",  "111110010111011001",  "111110010111011100",  "111110010111100000",  "111110010111100011",  "111110010111100110",  "111110010111101010",  "111110010111101101",  "111110010111110001",  "111110010111110101",  "111110010111111001",  "111110010111111100",  "111110011000000000",  "111110011000000100",  "111110011000001000",  "111110011000001100",  "111110011000010000",  "111110011000010101",  "111110011000011001",  "111110011000011101",  "111110011000100010",  "111110011000100110",  "111110011000101011",  "111110011000101111",  "111110011000110100",  "111110011000111000",  "111110011000111101",  "111110011001000010",  "111110011001000111",  "111110011001001100",  "111110011001010001",  "111110011001010110",  "111110011001011011",  "111110011001100001",  "111110011001100110",  "111110011001101011",  "111110011001110001",  "111110011001110110",  "111110011001111100",  "111110011010000001",  "111110011010000111",  "111110011010001101",  "111110011010010011",  "111110011010011000",  "111110011010011110",  "111110011010100100",  "111110011010101010",  "111110011010110001",  "111110011010110111",  "111110011010111101",  "111110011011000011",  "111110011011001010",  "111110011011010000",  "111110011011010111",  "111110011011011101",  "111110011011100100",  "111110011011101011",  "111110011011110001",  "111110011011111000",  "111110011011111111",  "111110011100000110",  "111110011100001101",  "111110011100010100",  "111110011100011011",  "111110011100100010",  "111110011100101010",  "111110011100110001",  "111110011100111000",  "111110011101000000",  "111110011101000111",  "111110011101001111",  "111110011101010111",  "111110011101011110",  "111110011101100110",  "111110011101101110",  "111110011101110110",  "111110011101111110",  "111110011110000110",  "111110011110001110",  "111110011110010110",  "111110011110011110",  "111110011110100111",  "111110011110101111",  "111110011110110111",  "111110011111000000",  "111110011111001000",  "111110011111010001",  "111110011111011010",  "111110011111100010",  "111110011111101011",  "111110011111110100",  "111110011111111101",  "111110100000000110",  "111110100000001111",  "111110100000011000",  "111110100000100001",  "111110100000101010",  "111110100000110100",  "111110100000111101",  "111110100001000110",  "111110100001010000",  "111110100001011001",  "111110100001100011",  "111110100001101100",  "111110100001110110",  "111110100010000000",  "111110100010001010",  "111110100010010100",  "111110100010011110",  "111110100010101000",  "111110100010110010",  "111110100010111100",  "111110100011000110",  "111110100011010000",  "111110100011011011",  "111110100011100101",  "111110100011101111",  "111110100011111010",  "111110100100000100",  "111110100100001111",  "111110100100011010",  "111110100100100100",  "111110100100101111",  "111110100100111010",  "111110100101000101",  "111110100101010000",  "111110100101011011",  "111110100101100110",  "111110100101110001",  "111110100101111101",  "111110100110001000",  "111110100110010011",  "111110100110011110",  "111110100110101010",  "111110100110110101",  "111110100111000001",  "111110100111001101",  "111110100111011000",  "111110100111100100",  "111110100111110000",  "111110100111111100",  "111110101000001000",  "111110101000010100",  "111110101000100000",  "111110101000101100",  "111110101000111000",  "111110101001000100",  "111110101001010000",  "111110101001011101",  "111110101001101001",  "111110101001110110",  "111110101010000010",  "111110101010001111",  "111110101010011011",  "111110101010101000",  "111110101010110101",  "111110101011000001",  "111110101011001110",  "111110101011011011",  "111110101011101000",  "111110101011110101",  "111110101100000010",  "111110101100001111",  "111110101100011101",  "111110101100101010",  "111110101100110111",  "111110101101000100",  "111110101101010010",  "111110101101011111",  "111110101101101101",  "111110101101111010",  "111110101110001000",  "111110101110010110",  "111110101110100100",  "111110101110110001",  "111110101110111111",  "111110101111001101",  "111110101111011011",  "111110101111101001",  "111110101111110111",  "111110110000000101",  "111110110000010011",  "111110110000100010",  "111110110000110000",  "111110110000111110",  "111110110001001101",  "111110110001011011",  "111110110001101010",  "111110110001111000",  "111110110010000111",  "111110110010010110",  "111110110010100100",  "111110110010110011",  "111110110011000010",  "111110110011010001",  "111110110011100000",  "111110110011101111",  "111110110011111110",  "111110110100001101",  "111110110100011100",  "111110110100101011",  "111110110100111010",  "111110110101001010",  "111110110101011001",  "111110110101101001",  "111110110101111000",  "111110110110001000",  "111110110110010111",  "111110110110100111",  "111110110110110110",  "111110110111000110",  "111110110111010110",  "111110110111100110",  "111110110111110110",  "111110111000000101",  "111110111000010101",  "111110111000100101",  "111110111000110110",  "111110111001000110",  "111110111001010110",  "111110111001100110",  "111110111001110110",  "111110111010000111",  "111110111010010111",  "111110111010101000",  "111110111010111000",  "111110111011001000",  "111110111011011001",  "111110111011101010",  "111110111011111010",  "111110111100001011",  "111110111100011100",  "111110111100101101",  "111110111100111110",  "111110111101001110",  "111110111101011111",  "111110111101110000",  "111110111110000001",  "111110111110010011",  "111110111110100100",  "111110111110110101",  "111110111111000110",  "111110111111010111",  "111110111111101001",  "111110111111111010",  "111111000000001100",  "111111000000011101",  "111111000000101111",  "111111000001000000",  "111111000001010010",  "111111000001100011",  "111111000001110101",  "111111000010000111",  "111111000010011001",  "111111000010101011",  "111111000010111100",  "111111000011001110",  "111111000011100000",  "111111000011110010",  "111111000100000101",  "111111000100010111",  "111111000100101001",  "111111000100111011",  "111111000101001101",  "111111000101100000",  "111111000101110010",  "111111000110000100",  "111111000110010111",  "111111000110101001",  "111111000110111100",  "111111000111001110",  "111111000111100001",  "111111000111110011",  "111111001000000110",  "111111001000011001",  "111111001000101100",  "111111001000111110",  "111111001001010001",  "111111001001100100",  "111111001001110111",  "111111001010001010",  "111111001010011101",  "111111001010110000",  "111111001011000011",  "111111001011010110",  "111111001011101010",  "111111001011111101",  "111111001100010000",  "111111001100100011",  "111111001100110111",  "111111001101001010",  "111111001101011101",  "111111001101110001",  "111111001110000100",  "111111001110011000",  "111111001110101011",  "111111001110111111",  "111111001111010011",  "111111001111100110",  "111111001111111010",  "111111010000001110",  "111111010000100010",  "111111010000110110",  "111111010001001001",  "111111010001011101",  "111111010001110001",  "111111010010000101",  "111111010010011001",  "111111010010101101",  "111111010011000001",  "111111010011010110",  "111111010011101010",  "111111010011111110",  "111111010100010010",  "111111010100100111",  "111111010100111011",  "111111010101001111",  "111111010101100100",  "111111010101111000",  "111111010110001100",  "111111010110100001",  "111111010110110101",  "111111010111001010",  "111111010111011111",  "111111010111110011",  "111111011000001000",  "111111011000011101",  "111111011000110001",  "111111011001000110",  "111111011001011011",  "111111011001110000",  "111111011010000101",  "111111011010011001",  "111111011010101110",  "111111011011000011",  "111111011011011000",  "111111011011101101",  "111111011100000010",  "111111011100010111",  "111111011100101101",  "111111011101000010",  "111111011101010111",  "111111011101101100",  "111111011110000001",  "111111011110010111",  "111111011110101100",  "111111011111000001",  "111111011111010111",  "111111011111101100",  "111111100000000001",  "111111100000010111",  "111111100000101100",  "111111100001000010",  "111111100001010111",  "111111100001101101",  "111111100010000011",  "111111100010011000",  "111111100010101110",  "111111100011000011",  "111111100011011001",  "111111100011101111",  "111111100100000101",  "111111100100011010",  "111111100100110000",  "111111100101000110",  "111111100101011100",  "111111100101110010",  "111111100110001000",  "111111100110011110",  "111111100110110100",  "111111100111001010",  "111111100111100000",  "111111100111110110",  "111111101000001100",  "111111101000100010",  "111111101000111000",  "111111101001001110",  "111111101001100100",  "111111101001111010",  "111111101010010001",  "111111101010100111",  "111111101010111101",  "111111101011010011",  "111111101011101010",  "111111101100000000",  "111111101100010110",  "111111101100101101",  "111111101101000011",  "111111101101011010",  "111111101101110000",  "111111101110000110",  "111111101110011101",  "111111101110110011",  "111111101111001010",  "111111101111100000",  "111111101111110111",  "111111110000001110",  "111111110000100100",  "111111110000111011",  "111111110001010001",  "111111110001101000",  "111111110001111111",  "111111110010010110",  "111111110010101100",  "111111110011000011",  "111111110011011010",  "111111110011110000",  "111111110100000111",  "111111110100011110",  "111111110100110101",  "111111110101001100",  "111111110101100011",  "111111110101111001",  "111111110110010000",  "111111110110100111",  "111111110110111110",  "111111110111010101",  "111111110111101100",  "111111111000000011",  "111111111000011010",  "111111111000110001",  "111111111001001000",  "111111111001011111",  "111111111001110110",  "111111111010001101",  "111111111010100100",  "111111111010111011",  "111111111011010010",  "111111111011101010",  "111111111100000001",  "111111111100011000",  "111111111100101111",  "111111111101000110",  "111111111101011101",  "111111111101110101",  "111111111110001100",  "111111111110100011",  "111111111110111010",  "111111111111010001",  "111111111111101001"),("000000000000000000",  "000000000000010111",  "000000000000101111",  "000000000001000110",  "000000000001011101",  "000000000001110100",  "000000000010001100",  "000000000010100011",  "000000000010111010",  "000000000011010010",  "000000000011101001",  "000000000100000001",  "000000000100011000",  "000000000100101111",  "000000000101000111",  "000000000101011110",  "000000000101110110",  "000000000110001101",  "000000000110100100",  "000000000110111100",  "000000000111010011",  "000000000111101011",  "000000001000000010",  "000000001000011010",  "000000001000110001",  "000000001001001001",  "000000001001100000",  "000000001001111000",  "000000001010001111",  "000000001010100111",  "000000001010111110",  "000000001011010110",  "000000001011101101",  "000000001100000101",  "000000001100011100",  "000000001100110100",  "000000001101001011",  "000000001101100011",  "000000001101111010",  "000000001110010010",  "000000001110101001",  "000000001111000001",  "000000001111011000",  "000000001111110000",  "000000010000000111",  "000000010000011111",  "000000010000110110",  "000000010001001110",  "000000010001100101",  "000000010001111101",  "000000010010010101",  "000000010010101100",  "000000010011000100",  "000000010011011011",  "000000010011110011",  "000000010100001010",  "000000010100100010",  "000000010100111001",  "000000010101010001",  "000000010101101000",  "000000010110000000",  "000000010110010111",  "000000010110101111",  "000000010111000111",  "000000010111011110",  "000000010111110110",  "000000011000001101",  "000000011000100101",  "000000011000111100",  "000000011001010100",  "000000011001101011",  "000000011010000011",  "000000011010011010",  "000000011010110010",  "000000011011001001",  "000000011011100001",  "000000011011111000",  "000000011100001111",  "000000011100100111",  "000000011100111110",  "000000011101010110",  "000000011101101101",  "000000011110000101",  "000000011110011100",  "000000011110110100",  "000000011111001011",  "000000011111100010",  "000000011111111010",  "000000100000010001",  "000000100000101000",  "000000100001000000",  "000000100001010111",  "000000100001101111",  "000000100010000110",  "000000100010011101",  "000000100010110101",  "000000100011001100",  "000000100011100011",  "000000100011111010",  "000000100100010010",  "000000100100101001",  "000000100101000000",  "000000100101011000",  "000000100101101111",  "000000100110000110",  "000000100110011101",  "000000100110110100",  "000000100111001100",  "000000100111100011",  "000000100111111010",  "000000101000010001",  "000000101000101000",  "000000101000111111",  "000000101001010110",  "000000101001101101",  "000000101010000101",  "000000101010011100",  "000000101010110011",  "000000101011001010",  "000000101011100001",  "000000101011111000",  "000000101100001111",  "000000101100100110",  "000000101100111101",  "000000101101010100",  "000000101101101011",  "000000101110000001",  "000000101110011000",  "000000101110101111",  "000000101111000110",  "000000101111011101",  "000000101111110100",  "000000110000001010",  "000000110000100001",  "000000110000111000",  "000000110001001111",  "000000110001100110",  "000000110001111100",  "000000110010010011",  "000000110010101010",  "000000110011000000",  "000000110011010111",  "000000110011101101",  "000000110100000100",  "000000110100011011",  "000000110100110001",  "000000110101001000",  "000000110101011110",  "000000110101110101",  "000000110110001011",  "000000110110100010",  "000000110110111000",  "000000110111001110",  "000000110111100101",  "000000110111111011",  "000000111000010001",  "000000111000101000",  "000000111000111110",  "000000111001010100",  "000000111001101011",  "000000111010000001",  "000000111010010111",  "000000111010101101",  "000000111011000011",  "000000111011011001",  "000000111011101111",  "000000111100000101",  "000000111100011011",  "000000111100110001",  "000000111101000111",  "000000111101011101",  "000000111101110011",  "000000111110001001",  "000000111110011111",  "000000111110110101",  "000000111111001011",  "000000111111100001",  "000000111111110110",  "000001000000001100",  "000001000000100010",  "000001000000110111",  "000001000001001101",  "000001000001100011",  "000001000001111000",  "000001000010001110",  "000001000010100011",  "000001000010111001",  "000001000011001110",  "000001000011100100",  "000001000011111001",  "000001000100001111",  "000001000100100100",  "000001000100111001",  "000001000101001110",  "000001000101100100",  "000001000101111001",  "000001000110001110",  "000001000110100011",  "000001000110111000",  "000001000111001101",  "000001000111100011",  "000001000111111000",  "000001001000001101",  "000001001000100010",  "000001001000110110",  "000001001001001011",  "000001001001100000",  "000001001001110101",  "000001001010001010",  "000001001010011111",  "000001001010110011",  "000001001011001000",  "000001001011011101",  "000001001011110001",  "000001001100000110",  "000001001100011010",  "000001001100101111",  "000001001101000011",  "000001001101011000",  "000001001101101100",  "000001001110000000",  "000001001110010101",  "000001001110101001",  "000001001110111101",  "000001001111010010",  "000001001111100110",  "000001001111111010",  "000001010000001110",  "000001010000100010",  "000001010000110110",  "000001010001001010",  "000001010001011110",  "000001010001110010",  "000001010010000110",  "000001010010011001",  "000001010010101101",  "000001010011000001",  "000001010011010101",  "000001010011101000",  "000001010011111100",  "000001010100001111",  "000001010100100011",  "000001010100110110",  "000001010101001010",  "000001010101011101",  "000001010101110001",  "000001010110000100",  "000001010110010111",  "000001010110101010",  "000001010110111110",  "000001010111010001",  "000001010111100100",  "000001010111110111",  "000001011000001010",  "000001011000011101",  "000001011000110000",  "000001011001000011",  "000001011001010110",  "000001011001101000",  "000001011001111011",  "000001011010001110",  "000001011010100000",  "000001011010110011",  "000001011011000110",  "000001011011011000",  "000001011011101011",  "000001011011111101",  "000001011100001111",  "000001011100100010",  "000001011100110100",  "000001011101000110",  "000001011101011000",  "000001011101101011",  "000001011101111101",  "000001011110001111",  "000001011110100001",  "000001011110110011",  "000001011111000101",  "000001011111010110",  "000001011111101000",  "000001011111111010",  "000001100000001100",  "000001100000011101",  "000001100000101111",  "000001100001000001",  "000001100001010010",  "000001100001100100",  "000001100001110101",  "000001100010000110",  "000001100010011000",  "000001100010101001",  "000001100010111010",  "000001100011001011",  "000001100011011100",  "000001100011101101",  "000001100011111110",  "000001100100001111",  "000001100100100000",  "000001100100110001",  "000001100101000010",  "000001100101010011",  "000001100101100011",  "000001100101110100",  "000001100110000100",  "000001100110010101",  "000001100110100101",  "000001100110110110",  "000001100111000110",  "000001100111010110",  "000001100111100111",  "000001100111110111",  "000001101000000111",  "000001101000010111",  "000001101000100111",  "000001101000110111",  "000001101001000111",  "000001101001010111",  "000001101001100111",  "000001101001110110",  "000001101010000110",  "000001101010010110",  "000001101010100101",  "000001101010110101",  "000001101011000100",  "000001101011010100",  "000001101011100011",  "000001101011110010",  "000001101100000010",  "000001101100010001",  "000001101100100000",  "000001101100101111",  "000001101100111110",  "000001101101001101",  "000001101101011100",  "000001101101101011",  "000001101101111001",  "000001101110001000",  "000001101110010111",  "000001101110100101",  "000001101110110100",  "000001101111000010",  "000001101111010001",  "000001101111011111",  "000001101111101101",  "000001101111111100",  "000001110000001010",  "000001110000011000",  "000001110000100110",  "000001110000110100",  "000001110001000010",  "000001110001010000",  "000001110001011110",  "000001110001101011",  "000001110001111001",  "000001110010000111",  "000001110010010100",  "000001110010100010",  "000001110010101111",  "000001110010111100",  "000001110011001010",  "000001110011010111",  "000001110011100100",  "000001110011110001",  "000001110011111110",  "000001110100001011",  "000001110100011000",  "000001110100100101",  "000001110100110010",  "000001110100111111",  "000001110101001011",  "000001110101011000",  "000001110101100100",  "000001110101110001",  "000001110101111101",  "000001110110001010",  "000001110110010110",  "000001110110100010",  "000001110110101110",  "000001110110111010",  "000001110111000110",  "000001110111010010",  "000001110111011110",  "000001110111101010",  "000001110111110110",  "000001111000000010",  "000001111000001101",  "000001111000011001",  "000001111000100100",  "000001111000110000",  "000001111000111011",  "000001111001000110",  "000001111001010001",  "000001111001011101",  "000001111001101000",  "000001111001110011",  "000001111001111110",  "000001111010001000",  "000001111010010011",  "000001111010011110",  "000001111010101001",  "000001111010110011",  "000001111010111110",  "000001111011001000",  "000001111011010011",  "000001111011011101",  "000001111011100111",  "000001111011110001",  "000001111011111100",  "000001111100000110",  "000001111100010000",  "000001111100011001",  "000001111100100011",  "000001111100101101",  "000001111100110111",  "000001111101000000",  "000001111101001010",  "000001111101010011",  "000001111101011101",  "000001111101100110",  "000001111101101111",  "000001111101111001",  "000001111110000010",  "000001111110001011",  "000001111110010100",  "000001111110011101",  "000001111110100110",  "000001111110101110",  "000001111110110111",  "000001111111000000",  "000001111111001000",  "000001111111010001",  "000001111111011001",  "000001111111100001",  "000001111111101010",  "000001111111110010",  "000001111111111010",  "000010000000000010",  "000010000000001010",  "000010000000010010",  "000010000000011010",  "000010000000100001",  "000010000000101001",  "000010000000110001",  "000010000000111000",  "000010000001000000",  "000010000001000111",  "000010000001001110",  "000010000001010101",  "000010000001011101",  "000010000001100100",  "000010000001101011",  "000010000001110010",  "000010000001111000",  "000010000001111111",  "000010000010000110",  "000010000010001101",  "000010000010010011",  "000010000010011010",  "000010000010100000",  "000010000010100110",  "000010000010101101",  "000010000010110011",  "000010000010111001",  "000010000010111111",  "000010000011000101",  "000010000011001011",  "000010000011010000",  "000010000011010110",  "000010000011011100",  "000010000011100001",  "000010000011100111",  "000010000011101100",  "000010000011110010",  "000010000011110111",  "000010000011111100",  "000010000100000001",  "000010000100000110",  "000010000100001011",  "000010000100010000",  "000010000100010101",  "000010000100011001",  "000010000100011110",  "000010000100100011",  "000010000100100111",  "000010000100101100",  "000010000100110000",  "000010000100110100",  "000010000100111000",  "000010000100111100",  "000010000101000000",  "000010000101000100",  "000010000101001000",  "000010000101001100",  "000010000101010000",  "000010000101010011",  "000010000101010111",  "000010000101011010",  "000010000101011110",  "000010000101100001",  "000010000101100100",  "000010000101100111",  "000010000101101010",  "000010000101101101",  "000010000101110000",  "000010000101110011",  "000010000101110110",  "000010000101111001",  "000010000101111011",  "000010000101111110",  "000010000110000000",  "000010000110000010",  "000010000110000101",  "000010000110000111",  "000010000110001001",  "000010000110001011",  "000010000110001101",  "000010000110001111",  "000010000110010001",  "000010000110010010",  "000010000110010100",  "000010000110010110",  "000010000110010111",  "000010000110011000",  "000010000110011010",  "000010000110011011",  "000010000110011100",  "000010000110011101",  "000010000110011110",  "000010000110011111",  "000010000110100000",  "000010000110100001",  "000010000110100001",  "000010000110100010",  "000010000110100010",  "000010000110100011",  "000010000110100011",  "000010000110100011",  "000010000110100100",  "000010000110100100",  "000010000110100100",  "000010000110100100",  "000010000110100011",  "000010000110100011",  "000010000110100011",  "000010000110100011",  "000010000110100010",  "000010000110100010",  "000010000110100001",  "000010000110100000",  "000010000110011111",  "000010000110011111",  "000010000110011110",  "000010000110011101",  "000010000110011011",  "000010000110011010",  "000010000110011001",  "000010000110011000",  "000010000110010110",  "000010000110010101",  "000010000110010011",  "000010000110010001",  "000010000110001111",  "000010000110001110",  "000010000110001100",  "000010000110001010",  "000010000110000111",  "000010000110000101",  "000010000110000011",  "000010000110000001",  "000010000101111110",  "000010000101111100",  "000010000101111001",  "000010000101110110",  "000010000101110100",  "000010000101110001",  "000010000101101110",  "000010000101101011",  "000010000101101000",  "000010000101100101",  "000010000101100001",  "000010000101011110",  "000010000101011011",  "000010000101010111",  "000010000101010011",  "000010000101010000",  "000010000101001100",  "000010000101001000",  "000010000101000100",  "000010000101000000",  "000010000100111100",  "000010000100111000",  "000010000100110100",  "000010000100101111",  "000010000100101011",  "000010000100100111",  "000010000100100010",  "000010000100011101",  "000010000100011001",  "000010000100010100",  "000010000100001111",  "000010000100001010",  "000010000100000101",  "000010000100000000",  "000010000011111010",  "000010000011110101",  "000010000011110000",  "000010000011101010",  "000010000011100101",  "000010000011011111",  "000010000011011001",  "000010000011010011",  "000010000011001110",  "000010000011001000",  "000010000011000010",  "000010000010111011",  "000010000010110101",  "000010000010101111",  "000010000010101000",  "000010000010100010",  "000010000010011011",  "000010000010010101",  "000010000010001110",  "000010000010000111",  "000010000010000000",  "000010000001111001",  "000010000001110010",  "000010000001101011",  "000010000001100100",  "000010000001011101",  "000010000001010101",  "000010000001001110",  "000010000001000110",  "000010000000111111",  "000010000000110111",  "000010000000101111",  "000010000000100111",  "000010000000100000",  "000010000000010111",  "000010000000001111",  "000010000000000111",  "000001111111111111",  "000001111111110111",  "000001111111101110",  "000001111111100110",  "000001111111011101",  "000001111111010100",  "000001111111001100",  "000001111111000011",  "000001111110111010",  "000001111110110001",  "000001111110101000",  "000001111110011111",  "000001111110010101",  "000001111110001100",  "000001111110000011",  "000001111101111001",  "000001111101110000",  "000001111101100110",  "000001111101011100",  "000001111101010010",  "000001111101001000",  "000001111100111110",  "000001111100110100",  "000001111100101010",  "000001111100100000",  "000001111100010110",  "000001111100001011",  "000001111100000001",  "000001111011110110",  "000001111011101100",  "000001111011100001",  "000001111011010110",  "000001111011001011",  "000001111011000000",  "000001111010110101",  "000001111010101010",  "000001111010011111",  "000001111010010100",  "000001111010001001",  "000001111001111101",  "000001111001110010",  "000001111001100110",  "000001111001011010",  "000001111001001111",  "000001111001000011",  "000001111000110111",  "000001111000101011",  "000001111000011111",  "000001111000010011",  "000001111000000111",  "000001110111111010",  "000001110111101110",  "000001110111100010",  "000001110111010101",  "000001110111001000",  "000001110110111100",  "000001110110101111",  "000001110110100010",  "000001110110010101",  "000001110110001000",  "000001110101111011",  "000001110101101110",  "000001110101100001",  "000001110101010011",  "000001110101000110",  "000001110100111001",  "000001110100101011",  "000001110100011101",  "000001110100010000",  "000001110100000010",  "000001110011110100",  "000001110011100110",  "000001110011011000",  "000001110011001010",  "000001110010111100",  "000001110010101110",  "000001110010011111",  "000001110010010001",  "000001110010000011",  "000001110001110100",  "000001110001100101",  "000001110001010111",  "000001110001001000",  "000001110000111001",  "000001110000101010",  "000001110000011011",  "000001110000001100",  "000001101111111101",  "000001101111101110",  "000001101111011110",  "000001101111001111",  "000001101111000000",  "000001101110110000",  "000001101110100000",  "000001101110010001",  "000001101110000001",  "000001101101110001",  "000001101101100001",  "000001101101010001",  "000001101101000001",  "000001101100110001",  "000001101100100001",  "000001101100010001",  "000001101100000000",  "000001101011110000",  "000001101011100000",  "000001101011001111",  "000001101010111110",  "000001101010101110",  "000001101010011101",  "000001101010001100",  "000001101001111011",  "000001101001101010",  "000001101001011001",  "000001101001001000",  "000001101000110111",  "000001101000100101",  "000001101000010100",  "000001101000000010",  "000001100111110001",  "000001100111011111",  "000001100111001110",  "000001100110111100",  "000001100110101010",  "000001100110011000",  "000001100110000110",  "000001100101110100",  "000001100101100010",  "000001100101010000",  "000001100100111110",  "000001100100101100",  "000001100100011001",  "000001100100000111",  "000001100011110100",  "000001100011100010",  "000001100011001111",  "000001100010111100",  "000001100010101010",  "000001100010010111",  "000001100010000100",  "000001100001110001",  "000001100001011110",  "000001100001001011",  "000001100000111000",  "000001100000100100",  "000001100000010001",  "000001011111111110",  "000001011111101010",  "000001011111010111",  "000001011111000011",  "000001011110101111",  "000001011110011011",  "000001011110001000",  "000001011101110100",  "000001011101100000",  "000001011101001100",  "000001011100111000",  "000001011100100100",  "000001011100001111",  "000001011011111011",  "000001011011100111",  "000001011011010010",  "000001011010111110",  "000001011010101001",  "000001011010010101",  "000001011010000000",  "000001011001101011",  "000001011001010111",  "000001011001000010",  "000001011000101101",  "000001011000011000",  "000001011000000011",  "000001010111101110",  "000001010111011000",  "000001010111000011",  "000001010110101110",  "000001010110011000",  "000001010110000011",  "000001010101101110",  "000001010101011000",  "000001010101000010",  "000001010100101101",  "000001010100010111",  "000001010100000001",  "000001010011101011",  "000001010011010101",  "000001010010111111",  "000001010010101001",  "000001010010010011",  "000001010001111101",  "000001010001100111",  "000001010001010000",  "000001010000111010",  "000001010000100011",  "000001010000001101",  "000001001111110110",  "000001001111100000",  "000001001111001001",  "000001001110110010",  "000001001110011100",  "000001001110000101",  "000001001101101110",  "000001001101010111",  "000001001101000000",  "000001001100101001",  "000001001100010010",  "000001001011111010",  "000001001011100011",  "000001001011001100",  "000001001010110100",  "000001001010011101",  "000001001010000101",  "000001001001101110",  "000001001001010110",  "000001001000111111",  "000001001000100111",  "000001001000001111",  "000001000111110111",  "000001000111011111",  "000001000111000111",  "000001000110101111",  "000001000110010111",  "000001000101111111",  "000001000101100111",  "000001000101001111",  "000001000100110111",  "000001000100011110",  "000001000100000110",  "000001000011101101",  "000001000011010101",  "000001000010111100",  "000001000010100100",  "000001000010001011",  "000001000001110010",  "000001000001011010",  "000001000001000001",  "000001000000101000",  "000001000000001111",  "000000111111110110",  "000000111111011101",  "000000111111000100",  "000000111110101011",  "000000111110010010",  "000000111101111000",  "000000111101011111",  "000000111101000110",  "000000111100101100",  "000000111100010011",  "000000111011111001",  "000000111011100000",  "000000111011000110",  "000000111010101101",  "000000111010010011",  "000000111001111001",  "000000111001100000",  "000000111001000110",  "000000111000101100",  "000000111000010010",  "000000110111111000",  "000000110111011110",  "000000110111000100",  "000000110110101010",  "000000110110010000",  "000000110101110101",  "000000110101011011",  "000000110101000001",  "000000110100100110",  "000000110100001100",  "000000110011110010",  "000000110011010111",  "000000110010111101",  "000000110010100010",  "000000110010000111",  "000000110001101101",  "000000110001010010",  "000000110000110111",  "000000110000011101",  "000000110000000010",  "000000101111100111",  "000000101111001100",  "000000101110110001",  "000000101110010110",  "000000101101111011",  "000000101101100000",  "000000101101000101",  "000000101100101001",  "000000101100001110",  "000000101011110011",  "000000101011011000",  "000000101010111100",  "000000101010100001",  "000000101010000101",  "000000101001101010",  "000000101001001111",  "000000101000110011",  "000000101000010111",  "000000100111111100",  "000000100111100000",  "000000100111000100",  "000000100110101001",  "000000100110001101",  "000000100101110001",  "000000100101010101",  "000000100100111001",  "000000100100011101",  "000000100100000001",  "000000100011100101",  "000000100011001001",  "000000100010101101",  "000000100010010001",  "000000100001110101",  "000000100001011001",  "000000100000111101",  "000000100000100000",  "000000100000000100",  "000000011111101000",  "000000011111001011",  "000000011110101111",  "000000011110010011",  "000000011101110110",  "000000011101011010",  "000000011100111101",  "000000011100100001",  "000000011100000100",  "000000011011100111",  "000000011011001011",  "000000011010101110",  "000000011010010001",  "000000011001110100",  "000000011001011000",  "000000011000111011",  "000000011000011110",  "000000011000000001",  "000000010111100100",  "000000010111000111",  "000000010110101010",  "000000010110001101",  "000000010101110000",  "000000010101010011",  "000000010100110110",  "000000010100011001",  "000000010011111100",  "000000010011011111",  "000000010011000010",  "000000010010100100",  "000000010010000111",  "000000010001101010",  "000000010001001101",  "000000010000101111",  "000000010000010010",  "000000001111110100",  "000000001111010111",  "000000001110111010",  "000000001110011100",  "000000001101111111",  "000000001101100001",  "000000001101000100",  "000000001100100110",  "000000001100001000",  "000000001011101011",  "000000001011001101",  "000000001010110000",  "000000001010010010",  "000000001001110100",  "000000001001010111",  "000000001000111001",  "000000001000011011",  "000000000111111101",  "000000000111011111",  "000000000111000010",  "000000000110100100",  "000000000110000110",  "000000000101101000",  "000000000101001010",  "000000000100101100",  "000000000100001110",  "000000000011110000",  "000000000011010010",  "000000000010110100",  "000000000010010110",  "000000000001111000",  "000000000001011010",  "000000000000111100",  "000000000000011110"),("000000000000000000",  "111111111111100010",  "111111111111000100",  "111111111110100110",  "111111111110000111",  "111111111101101001",  "111111111101001011",  "111111111100101101",  "111111111100001111",  "111111111011110000",  "111111111011010010",  "111111111010110100",  "111111111010010110",  "111111111001110111",  "111111111001011001",  "111111111000111011",  "111111111000011100",  "111111110111111110",  "111111110111100000",  "111111110111000001",  "111111110110100011",  "111111110110000100",  "111111110101100110",  "111111110101001000",  "111111110100101001",  "111111110100001011",  "111111110011101100",  "111111110011001110",  "111111110010101111",  "111111110010010001",  "111111110001110011",  "111111110001010100",  "111111110000110110",  "111111110000010111",  "111111101111111001",  "111111101111011010",  "111111101110111011",  "111111101110011101",  "111111101101111110",  "111111101101100000",  "111111101101000001",  "111111101100100011",  "111111101100000100",  "111111101011100110",  "111111101011000111",  "111111101010101001",  "111111101010001010",  "111111101001101011",  "111111101001001101",  "111111101000101110",  "111111101000010000",  "111111100111110001",  "111111100111010010",  "111111100110110100",  "111111100110010101",  "111111100101110111",  "111111100101011000",  "111111100100111001",  "111111100100011011",  "111111100011111100",  "111111100011011110",  "111111100010111111",  "111111100010100000",  "111111100010000010",  "111111100001100011",  "111111100001000101",  "111111100000100110",  "111111100000000111",  "111111011111101001",  "111111011111001010",  "111111011110101100",  "111111011110001101",  "111111011101101111",  "111111011101010000",  "111111011100110001",  "111111011100010011",  "111111011011110100",  "111111011011010110",  "111111011010110111",  "111111011010011001",  "111111011001111010",  "111111011001011011",  "111111011000111101",  "111111011000011110",  "111111011000000000",  "111111010111100001",  "111111010111000011",  "111111010110100100",  "111111010110000110",  "111111010101100111",  "111111010101001001",  "111111010100101011",  "111111010100001100",  "111111010011101110",  "111111010011001111",  "111111010010110001",  "111111010010010010",  "111111010001110100",  "111111010001010110",  "111111010000110111",  "111111010000011001",  "111111001111111010",  "111111001111011100",  "111111001110111110",  "111111001110100000",  "111111001110000001",  "111111001101100011",  "111111001101000101",  "111111001100100110",  "111111001100001000",  "111111001011101010",  "111111001011001100",  "111111001010101101",  "111111001010001111",  "111111001001110001",  "111111001001010011",  "111111001000110101",  "111111001000010111",  "111111000111111001",  "111111000111011010",  "111111000110111100",  "111111000110011110",  "111111000110000000",  "111111000101100010",  "111111000101000100",  "111111000100100110",  "111111000100001000",  "111111000011101010",  "111111000011001100",  "111111000010101111",  "111111000010010001",  "111111000001110011",  "111111000001010101",  "111111000000110111",  "111111000000011001",  "111110111111111100",  "111110111111011110",  "111110111111000000",  "111110111110100010",  "111110111110000101",  "111110111101100111",  "111110111101001001",  "111110111100101100",  "111110111100001110",  "111110111011110000",  "111110111011010011",  "111110111010110101",  "111110111010011000",  "111110111001111010",  "111110111001011101",  "111110111001000000",  "111110111000100010",  "111110111000000101",  "111110110111100111",  "111110110111001010",  "111110110110101101",  "111110110110010000",  "111110110101110010",  "111110110101010101",  "111110110100111000",  "111110110100011011",  "111110110011111110",  "111110110011100001",  "111110110011000100",  "111110110010100111",  "111110110010001010",  "111110110001101101",  "111110110001010000",  "111110110000110011",  "111110110000010110",  "111110101111111001",  "111110101111011100",  "111110101110111111",  "111110101110100011",  "111110101110000110",  "111110101101101001",  "111110101101001101",  "111110101100110000",  "111110101100010011",  "111110101011110111",  "111110101011011010",  "111110101010111110",  "111110101010100010",  "111110101010000101",  "111110101001101001",  "111110101001001100",  "111110101000110000",  "111110101000010100",  "111110100111111000",  "111110100111011011",  "111110100110111111",  "111110100110100011",  "111110100110000111",  "111110100101101011",  "111110100101001111",  "111110100100110011",  "111110100100010111",  "111110100011111011",  "111110100011100000",  "111110100011000100",  "111110100010101000",  "111110100010001100",  "111110100001110001",  "111110100001010101",  "111110100000111001",  "111110100000011110",  "111110100000000010",  "111110011111100111",  "111110011111001011",  "111110011110110000",  "111110011110010101",  "111110011101111001",  "111110011101011110",  "111110011101000011",  "111110011100101000",  "111110011100001101",  "111110011011110010",  "111110011011010111",  "111110011010111100",  "111110011010100001",  "111110011010000110",  "111110011001101011",  "111110011001010000",  "111110011000110101",  "111110011000011011",  "111110011000000000",  "111110010111100101",  "111110010111001011",  "111110010110110000",  "111110010110010110",  "111110010101111011",  "111110010101100001",  "111110010101000111",  "111110010100101100",  "111110010100010010",  "111110010011111000",  "111110010011011110",  "111110010011000100",  "111110010010101010",  "111110010010010000",  "111110010001110110",  "111110010001011100",  "111110010001000010",  "111110010000101001",  "111110010000001111",  "111110001111110101",  "111110001111011100",  "111110001111000010",  "111110001110101000",  "111110001110001111",  "111110001101110110",  "111110001101011100",  "111110001101000011",  "111110001100101010",  "111110001100010001",  "111110001011111000",  "111110001011011110",  "111110001011000101",  "111110001010101101",  "111110001010010100",  "111110001001111011",  "111110001001100010",  "111110001001001001",  "111110001000110001",  "111110001000011000",  "111110001000000000",  "111110000111100111",  "111110000111001111",  "111110000110110110",  "111110000110011110",  "111110000110000110",  "111110000101101101",  "111110000101010101",  "111110000100111101",  "111110000100100101",  "111110000100001101",  "111110000011110101",  "111110000011011110",  "111110000011000110",  "111110000010101110",  "111110000010010110",  "111110000001111111",  "111110000001100111",  "111110000001010000",  "111110000000111001",  "111110000000100001",  "111110000000001010",  "111101111111110011",  "111101111111011100",  "111101111111000101",  "111101111110101110",  "111101111110010111",  "111101111110000000",  "111101111101101001",  "111101111101010010",  "111101111100111011",  "111101111100100101",  "111101111100001110",  "111101111011111000",  "111101111011100001",  "111101111011001011",  "111101111010110101",  "111101111010011111",  "111101111010001000",  "111101111001110010",  "111101111001011100",  "111101111001000110",  "111101111000110000",  "111101111000011011",  "111101111000000101",  "111101110111101111",  "111101110111011010",  "111101110111000100",  "111101110110101111",  "111101110110011001",  "111101110110000100",  "111101110101101111",  "111101110101011010",  "111101110101000100",  "111101110100101111",  "111101110100011010",  "111101110100000110",  "111101110011110001",  "111101110011011100",  "111101110011000111",  "111101110010110011",  "111101110010011110",  "111101110010001010",  "111101110001110101",  "111101110001100001",  "111101110001001101",  "111101110000111001",  "111101110000100101",  "111101110000010001",  "111101101111111101",  "111101101111101001",  "111101101111010101",  "111101101111000001",  "111101101110101110",  "111101101110011010",  "111101101110000111",  "111101101101110011",  "111101101101100000",  "111101101101001101",  "111101101100111001",  "111101101100100110",  "111101101100010011",  "111101101100000000",  "111101101011101110",  "111101101011011011",  "111101101011001000",  "111101101010110110",  "111101101010100011",  "111101101010010001",  "111101101001111110",  "111101101001101100",  "111101101001011010",  "111101101001000111",  "111101101000110101",  "111101101000100011",  "111101101000010010",  "111101101000000000",  "111101100111101110",  "111101100111011100",  "111101100111001011",  "111101100110111001",  "111101100110101000",  "111101100110010111",  "111101100110000101",  "111101100101110100",  "111101100101100011",  "111101100101010010",  "111101100101000001",  "111101100100110000",  "111101100100100000",  "111101100100001111",  "111101100011111110",  "111101100011101110",  "111101100011011101",  "111101100011001101",  "111101100010111101",  "111101100010101101",  "111101100010011101",  "111101100010001101",  "111101100001111101",  "111101100001101101",  "111101100001011101",  "111101100001001110",  "111101100000111110",  "111101100000101111",  "111101100000011111",  "111101100000010000",  "111101100000000001",  "111101011111110010",  "111101011111100011",  "111101011111010100",  "111101011111000101",  "111101011110110110",  "111101011110100111",  "111101011110011001",  "111101011110001010",  "111101011101111100",  "111101011101101110",  "111101011101011111",  "111101011101010001",  "111101011101000011",  "111101011100110101",  "111101011100100111",  "111101011100011001",  "111101011100001100",  "111101011011111110",  "111101011011110001",  "111101011011100011",  "111101011011010110",  "111101011011001001",  "111101011010111100",  "111101011010101111",  "111101011010100010",  "111101011010010101",  "111101011010001000",  "111101011001111011",  "111101011001101111",  "111101011001100010",  "111101011001010110",  "111101011001001001",  "111101011000111101",  "111101011000110001",  "111101011000100101",  "111101011000011001",  "111101011000001101",  "111101011000000010",  "111101010111110110",  "111101010111101010",  "111101010111011111",  "111101010111010100",  "111101010111001000",  "111101010110111101",  "111101010110110010",  "111101010110100111",  "111101010110011100",  "111101010110010001",  "111101010110000111",  "111101010101111100",  "111101010101110010",  "111101010101100111",  "111101010101011101",  "111101010101010011",  "111101010101001001",  "111101010100111111",  "111101010100110101",  "111101010100101011",  "111101010100100001",  "111101010100010111",  "111101010100001110",  "111101010100000100",  "111101010011111011",  "111101010011110010",  "111101010011101001",  "111101010011100000",  "111101010011010111",  "111101010011001110",  "111101010011000101",  "111101010010111101",  "111101010010110100",  "111101010010101100",  "111101010010100011",  "111101010010011011",  "111101010010010011",  "111101010010001011",  "111101010010000011",  "111101010001111011",  "111101010001110011",  "111101010001101100",  "111101010001100100",  "111101010001011101",  "111101010001010101",  "111101010001001110",  "111101010001000111",  "111101010001000000",  "111101010000111001",  "111101010000110010",  "111101010000101011",  "111101010000100101",  "111101010000011110",  "111101010000011000",  "111101010000010001",  "111101010000001011",  "111101010000000101",  "111101001111111111",  "111101001111111001",  "111101001111110011",  "111101001111101110",  "111101001111101000",  "111101001111100011",  "111101001111011101",  "111101001111011000",  "111101001111010011",  "111101001111001110",  "111101001111001001",  "111101001111000100",  "111101001110111111",  "111101001110111010",  "111101001110110110",  "111101001110110001",  "111101001110101101",  "111101001110101001",  "111101001110100100",  "111101001110100000",  "111101001110011100",  "111101001110011001",  "111101001110010101",  "111101001110010001",  "111101001110001110",  "111101001110001010",  "111101001110000111",  "111101001110000100",  "111101001110000001",  "111101001101111110",  "111101001101111011",  "111101001101111000",  "111101001101110101",  "111101001101110011",  "111101001101110000",  "111101001101101110",  "111101001101101100",  "111101001101101001",  "111101001101100111",  "111101001101100101",  "111101001101100100",  "111101001101100010",  "111101001101100000",  "111101001101011111",  "111101001101011101",  "111101001101011100",  "111101001101011011",  "111101001101011010",  "111101001101011001",  "111101001101011000",  "111101001101010111",  "111101001101010111",  "111101001101010110",  "111101001101010110",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010110",  "111101001101010110",  "111101001101010111",  "111101001101010111",  "111101001101011000",  "111101001101011001",  "111101001101011010",  "111101001101011011",  "111101001101011100",  "111101001101011101",  "111101001101011111",  "111101001101100000",  "111101001101100010",  "111101001101100100",  "111101001101100101",  "111101001101100111",  "111101001101101001",  "111101001101101100",  "111101001101101110",  "111101001101110000",  "111101001101110011",  "111101001101110101",  "111101001101111000",  "111101001101111011",  "111101001101111110",  "111101001110000001",  "111101001110000100",  "111101001110000111",  "111101001110001011",  "111101001110001110",  "111101001110010010",  "111101001110010101",  "111101001110011001",  "111101001110011101",  "111101001110100001",  "111101001110100101",  "111101001110101001",  "111101001110101110",  "111101001110110010",  "111101001110110111",  "111101001110111100",  "111101001111000000",  "111101001111000101",  "111101001111001010",  "111101001111001111",  "111101001111010101",  "111101001111011010",  "111101001111011111",  "111101001111100101",  "111101001111101011",  "111101001111110000",  "111101001111110110",  "111101001111111100",  "111101010000000010",  "111101010000001001",  "111101010000001111",  "111101010000010101",  "111101010000011100",  "111101010000100011",  "111101010000101001",  "111101010000110000",  "111101010000110111",  "111101010000111110",  "111101010001000110",  "111101010001001101",  "111101010001010100",  "111101010001011100",  "111101010001100100",  "111101010001101011",  "111101010001110011",  "111101010001111011",  "111101010010000011",  "111101010010001011",  "111101010010010100",  "111101010010011100",  "111101010010100101",  "111101010010101101",  "111101010010110110",  "111101010010111111",  "111101010011001000",  "111101010011010001",  "111101010011011010",  "111101010011100100",  "111101010011101101",  "111101010011110110",  "111101010100000000",  "111101010100001010",  "111101010100010100",  "111101010100011110",  "111101010100101000",  "111101010100110010",  "111101010100111100",  "111101010101000111",  "111101010101010001",  "111101010101011100",  "111101010101100111",  "111101010101110001",  "111101010101111100",  "111101010110000111",  "111101010110010011",  "111101010110011110",  "111101010110101001",  "111101010110110101",  "111101010111000000",  "111101010111001100",  "111101010111011000",  "111101010111100100",  "111101010111110000",  "111101010111111100",  "111101011000001000",  "111101011000010101",  "111101011000100001",  "111101011000101110",  "111101011000111010",  "111101011001000111",  "111101011001010100",  "111101011001100001",  "111101011001101110",  "111101011001111100",  "111101011010001001",  "111101011010010110",  "111101011010100100",  "111101011010110010",  "111101011010111111",  "111101011011001101",  "111101011011011011",  "111101011011101001",  "111101011011111000",  "111101011100000110",  "111101011100010100",  "111101011100100011",  "111101011100110010",  "111101011101000000",  "111101011101001111",  "111101011101011110",  "111101011101101101",  "111101011101111101",  "111101011110001100",  "111101011110011011",  "111101011110101011",  "111101011110111010",  "111101011111001010",  "111101011111011010",  "111101011111101010",  "111101011111111010",  "111101100000001010",  "111101100000011010",  "111101100000101011",  "111101100000111011",  "111101100001001100",  "111101100001011101",  "111101100001101101",  "111101100001111110",  "111101100010001111",  "111101100010100000",  "111101100010110010",  "111101100011000011",  "111101100011010100",  "111101100011100110",  "111101100011111000",  "111101100100001001",  "111101100100011011",  "111101100100101101",  "111101100100111111",  "111101100101010001",  "111101100101100100",  "111101100101110110",  "111101100110001001",  "111101100110011011",  "111101100110101110",  "111101100111000001",  "111101100111010100",  "111101100111100111",  "111101100111111010",  "111101101000001101",  "111101101000100000",  "111101101000110100",  "111101101001000111",  "111101101001011011",  "111101101001101111",  "111101101010000010",  "111101101010010110",  "111101101010101010",  "111101101010111111",  "111101101011010011",  "111101101011100111",  "111101101011111100",  "111101101100010000",  "111101101100100101",  "111101101100111010",  "111101101101001110",  "111101101101100011",  "111101101101111000",  "111101101110001110",  "111101101110100011",  "111101101110111000",  "111101101111001110",  "111101101111100011",  "111101101111111001",  "111101110000001111",  "111101110000100101",  "111101110000111011",  "111101110001010001",  "111101110001100111",  "111101110001111101",  "111101110010010100",  "111101110010101010",  "111101110011000001",  "111101110011010111",  "111101110011101110",  "111101110100000101",  "111101110100011100",  "111101110100110011",  "111101110101001010",  "111101110101100010",  "111101110101111001",  "111101110110010001",  "111101110110101000",  "111101110111000000",  "111101110111011000",  "111101110111101111",  "111101111000000111",  "111101111000011111",  "111101111000111000",  "111101111001010000",  "111101111001101000",  "111101111010000001",  "111101111010011001",  "111101111010110010",  "111101111011001011",  "111101111011100100",  "111101111011111100",  "111101111100010110",  "111101111100101111",  "111101111101001000",  "111101111101100001",  "111101111101111011",  "111101111110010100",  "111101111110101110",  "111101111111000111",  "111101111111100001",  "111101111111111011",  "111110000000010101",  "111110000000101111",  "111110000001001001",  "111110000001100100",  "111110000001111110",  "111110000010011000",  "111110000010110011",  "111110000011001110",  "111110000011101000",  "111110000100000011",  "111110000100011110",  "111110000100111001",  "111110000101010100",  "111110000101101111",  "111110000110001011",  "111110000110100110",  "111110000111000010",  "111110000111011101",  "111110000111111001",  "111110001000010101",  "111110001000110000",  "111110001001001100",  "111110001001101000",  "111110001010000100",  "111110001010100001",  "111110001010111101",  "111110001011011001",  "111110001011110110",  "111110001100010010",  "111110001100101111",  "111110001101001100",  "111110001101101000",  "111110001110000101",  "111110001110100010",  "111110001110111111",  "111110001111011101",  "111110001111111010",  "111110010000010111",  "111110010000110101",  "111110010001010010",  "111110010001110000",  "111110010010001101",  "111110010010101011",  "111110010011001001",  "111110010011100111",  "111110010100000101",  "111110010100100011",  "111110010101000001",  "111110010101100000",  "111110010101111110",  "111110010110011100",  "111110010110111011",  "111110010111011010",  "111110010111111000",  "111110011000010111",  "111110011000110110",  "111110011001010101",  "111110011001110100",  "111110011010010011",  "111110011010110010",  "111110011011010010",  "111110011011110001",  "111110011100010000",  "111110011100110000",  "111110011101010000",  "111110011101101111",  "111110011110001111",  "111110011110101111",  "111110011111001111",  "111110011111101111",  "111110100000001111",  "111110100000101111",  "111110100001001111",  "111110100001110000",  "111110100010010000",  "111110100010110000",  "111110100011010001",  "111110100011110010",  "111110100100010010",  "111110100100110011",  "111110100101010100",  "111110100101110101",  "111110100110010110",  "111110100110110111",  "111110100111011000",  "111110100111111010",  "111110101000011011",  "111110101000111100",  "111110101001011110",  "111110101001111111",  "111110101010100001",  "111110101011000011",  "111110101011100100",  "111110101100000110",  "111110101100101000",  "111110101101001010",  "111110101101101100",  "111110101110001110",  "111110101110110001",  "111110101111010011",  "111110101111110101",  "111110110000011000",  "111110110000111010",  "111110110001011101",  "111110110001111111",  "111110110010100010",  "111110110011000101",  "111110110011101000",  "111110110100001011",  "111110110100101110",  "111110110101010001",  "111110110101110100",  "111110110110010111",  "111110110110111010",  "111110110111011101",  "111110111000000001",  "111110111000100100",  "111110111001001000",  "111110111001101011",  "111110111010001111",  "111110111010110011",  "111110111011010111",  "111110111011111010",  "111110111100011110",  "111110111101000010",  "111110111101100110",  "111110111110001011",  "111110111110101111",  "111110111111010011",  "111110111111110111",  "111111000000011100",  "111111000001000000",  "111111000001100101",  "111111000010001001",  "111111000010101110",  "111111000011010011",  "111111000011110111",  "111111000100011100",  "111111000101000001",  "111111000101100110",  "111111000110001011",  "111111000110110000",  "111111000111010101",  "111111000111111010",  "111111001000011111",  "111111001001000101",  "111111001001101010",  "111111001010001111",  "111111001010110101",  "111111001011011010",  "111111001100000000",  "111111001100100110",  "111111001101001011",  "111111001101110001",  "111111001110010111",  "111111001110111101",  "111111001111100011",  "111111010000001001",  "111111010000101111",  "111111010001010101",  "111111010001111011",  "111111010010100001",  "111111010011000111",  "111111010011101110",  "111111010100010100",  "111111010100111010",  "111111010101100001",  "111111010110000111",  "111111010110101110",  "111111010111010100",  "111111010111111011",  "111111011000100010",  "111111011001001001",  "111111011001101111",  "111111011010010110",  "111111011010111101",  "111111011011100100",  "111111011100001011",  "111111011100110010",  "111111011101011001",  "111111011110000000",  "111111011110101000",  "111111011111001111",  "111111011111110110",  "111111100000011110",  "111111100001000101",  "111111100001101100",  "111111100010010100",  "111111100010111011",  "111111100011100011",  "111111100100001011",  "111111100100110010",  "111111100101011010",  "111111100110000010",  "111111100110101001",  "111111100111010001",  "111111100111111001",  "111111101000100001",  "111111101001001001",  "111111101001110001",  "111111101010011001",  "111111101011000001",  "111111101011101001",  "111111101100010001",  "111111101100111001",  "111111101101100010",  "111111101110001010",  "111111101110110010",  "111111101111011011",  "111111110000000011",  "111111110000101011",  "111111110001010100",  "111111110001111100",  "111111110010100101",  "111111110011001110",  "111111110011110110",  "111111110100011111",  "111111110101000111",  "111111110101110000",  "111111110110011001",  "111111110111000010",  "111111110111101011",  "111111111000010011",  "111111111000111100",  "111111111001100101",  "111111111010001110",  "111111111010110111",  "111111111011100000",  "111111111100001001",  "111111111100110010",  "111111111101011011",  "111111111110000100",  "111111111110101110",  "111111111111010111"),("000000000000000000",  "000000000000101001",  "000000000001010011",  "000000000001111100",  "000000000010100101",  "000000000011001111",  "000000000011111000",  "000000000100100001",  "000000000101001011",  "000000000101110100",  "000000000110011110",  "000000000111000111",  "000000000111110001",  "000000001000011010",  "000000001001000100",  "000000001001101110",  "000000001010010111",  "000000001011000001",  "000000001011101011",  "000000001100010100",  "000000001100111110",  "000000001101101000",  "000000001110010001",  "000000001110111011",  "000000001111100101",  "000000010000001111",  "000000010000111001",  "000000010001100011",  "000000010010001100",  "000000010010110110",  "000000010011100000",  "000000010100001010",  "000000010100110100",  "000000010101011110",  "000000010110001000",  "000000010110110010",  "000000010111011100",  "000000011000000110",  "000000011000110000",  "000000011001011010",  "000000011010000100",  "000000011010101111",  "000000011011011001",  "000000011100000011",  "000000011100101101",  "000000011101010111",  "000000011110000001",  "000000011110101011",  "000000011111010110",  "000000100000000000",  "000000100000101010",  "000000100001010100",  "000000100001111110",  "000000100010101001",  "000000100011010011",  "000000100011111101",  "000000100100100111",  "000000100101010010",  "000000100101111100",  "000000100110100110",  "000000100111010000",  "000000100111111011",  "000000101000100101",  "000000101001001111",  "000000101001111010",  "000000101010100100",  "000000101011001110",  "000000101011111001",  "000000101100100011",  "000000101101001101",  "000000101101111000",  "000000101110100010",  "000000101111001100",  "000000101111110111",  "000000110000100001",  "000000110001001011",  "000000110001110110",  "000000110010100000",  "000000110011001010",  "000000110011110101",  "000000110100011111",  "000000110101001001",  "000000110101110100",  "000000110110011110",  "000000110111001000",  "000000110111110011",  "000000111000011101",  "000000111001000111",  "000000111001110010",  "000000111010011100",  "000000111011000110",  "000000111011110000",  "000000111100011011",  "000000111101000101",  "000000111101101111",  "000000111110011010",  "000000111111000100",  "000000111111101110",  "000001000000011000",  "000001000001000011",  "000001000001101101",  "000001000010010111",  "000001000011000001",  "000001000011101011",  "000001000100010110",  "000001000101000000",  "000001000101101010",  "000001000110010100",  "000001000110111110",  "000001000111101000",  "000001001000010011",  "000001001000111101",  "000001001001100111",  "000001001010010001",  "000001001010111011",  "000001001011100101",  "000001001100001111",  "000001001100111001",  "000001001101100011",  "000001001110001101",  "000001001110110111",  "000001001111100001",  "000001010000001011",  "000001010000110101",  "000001010001011111",  "000001010010001000",  "000001010010110010",  "000001010011011100",  "000001010100000110",  "000001010100110000",  "000001010101011010",  "000001010110000011",  "000001010110101101",  "000001010111010111",  "000001011000000000",  "000001011000101010",  "000001011001010100",  "000001011001111101",  "000001011010100111",  "000001011011010001",  "000001011011111010",  "000001011100100100",  "000001011101001101",  "000001011101110111",  "000001011110100000",  "000001011111001001",  "000001011111110011",  "000001100000011100",  "000001100001000101",  "000001100001101111",  "000001100010011000",  "000001100011000001",  "000001100011101010",  "000001100100010100",  "000001100100111101",  "000001100101100110",  "000001100110001111",  "000001100110111000",  "000001100111100001",  "000001101000001010",  "000001101000110011",  "000001101001011100",  "000001101010000101",  "000001101010101110",  "000001101011010111",  "000001101011111111",  "000001101100101000",  "000001101101010001",  "000001101101111001",  "000001101110100010",  "000001101111001011",  "000001101111110011",  "000001110000011100",  "000001110001000100",  "000001110001101101",  "000001110010010101",  "000001110010111110",  "000001110011100110",  "000001110100001110",  "000001110100110110",  "000001110101011111",  "000001110110000111",  "000001110110101111",  "000001110111010111",  "000001110111111111",  "000001111000100111",  "000001111001001111",  "000001111001110111",  "000001111010011111",  "000001111011000111",  "000001111011101110",  "000001111100010110",  "000001111100111110",  "000001111101100110",  "000001111110001101",  "000001111110110101",  "000001111111011100",  "000010000000000100",  "000010000000101011",  "000010000001010010",  "000010000001111010",  "000010000010100001",  "000010000011001000",  "000010000011101111",  "000010000100010110",  "000010000100111110",  "000010000101100101",  "000010000110001011",  "000010000110110010",  "000010000111011001",  "000010001000000000",  "000010001000100111",  "000010001001001101",  "000010001001110100",  "000010001010011011",  "000010001011000001",  "000010001011101000",  "000010001100001110",  "000010001100110100",  "000010001101011011",  "000010001110000001",  "000010001110100111",  "000010001111001101",  "000010001111110011",  "000010010000011001",  "000010010000111111",  "000010010001100101",  "000010010010001011",  "000010010010110001",  "000010010011010111",  "000010010011111100",  "000010010100100010",  "000010010101000111",  "000010010101101101",  "000010010110010010",  "000010010110111000",  "000010010111011101",  "000010011000000010",  "000010011000100111",  "000010011001001100",  "000010011001110001",  "000010011010010110",  "000010011010111011",  "000010011011100000",  "000010011100000101",  "000010011100101001",  "000010011101001110",  "000010011101110011",  "000010011110010111",  "000010011110111100",  "000010011111100000",  "000010100000000100",  "000010100000101000",  "000010100001001101",  "000010100001110001",  "000010100010010101",  "000010100010111001",  "000010100011011100",  "000010100100000000",  "000010100100100100",  "000010100101001000",  "000010100101101011",  "000010100110001111",  "000010100110110010",  "000010100111010101",  "000010100111111001",  "000010101000011100",  "000010101000111111",  "000010101001100010",  "000010101010000101",  "000010101010101000",  "000010101011001011",  "000010101011101101",  "000010101100010000",  "000010101100110011",  "000010101101010101",  "000010101101111000",  "000010101110011010",  "000010101110111100",  "000010101111011110",  "000010110000000001",  "000010110000100011",  "000010110001000101",  "000010110001100110",  "000010110010001000",  "000010110010101010",  "000010110011001100",  "000010110011101101",  "000010110100001111",  "000010110100110000",  "000010110101010001",  "000010110101110010",  "000010110110010100",  "000010110110110101",  "000010110111010110",  "000010110111110110",  "000010111000010111",  "000010111000111000",  "000010111001011001",  "000010111001111001",  "000010111010011001",  "000010111010111010",  "000010111011011010",  "000010111011111010",  "000010111100011010",  "000010111100111010",  "000010111101011010",  "000010111101111010",  "000010111110011010",  "000010111110111001",  "000010111111011001",  "000010111111111000",  "000011000000011000",  "000011000000110111",  "000011000001010110",  "000011000001110101",  "000011000010010100",  "000011000010110011",  "000011000011010010",  "000011000011110001",  "000011000100001111",  "000011000100101110",  "000011000101001100",  "000011000101101010",  "000011000110001001",  "000011000110100111",  "000011000111000101",  "000011000111100011",  "000011001000000001",  "000011001000011110",  "000011001000111100",  "000011001001011010",  "000011001001110111",  "000011001010010100",  "000011001010110010",  "000011001011001111",  "000011001011101100",  "000011001100001001",  "000011001100100110",  "000011001101000010",  "000011001101011111",  "000011001101111011",  "000011001110011000",  "000011001110110100",  "000011001111010000",  "000011001111101101",  "000011010000001001",  "000011010000100101",  "000011010001000000",  "000011010001011100",  "000011010001111000",  "000011010010010011",  "000011010010101111",  "000011010011001010",  "000011010011100101",  "000011010100000000",  "000011010100011011",  "000011010100110110",  "000011010101010001",  "000011010101101011",  "000011010110000110",  "000011010110100000",  "000011010110111011",  "000011010111010101",  "000011010111101111",  "000011011000001001",  "000011011000100011",  "000011011000111101",  "000011011001010110",  "000011011001110000",  "000011011010001001",  "000011011010100011",  "000011011010111100",  "000011011011010101",  "000011011011101110",  "000011011100000111",  "000011011100011111",  "000011011100111000",  "000011011101010001",  "000011011101101001",  "000011011110000001",  "000011011110011010",  "000011011110110010",  "000011011111001010",  "000011011111100001",  "000011011111111001",  "000011100000010001",  "000011100000101000",  "000011100001000000",  "000011100001010111",  "000011100001101110",  "000011100010000101",  "000011100010011100",  "000011100010110011",  "000011100011001001",  "000011100011100000",  "000011100011110110",  "000011100100001101",  "000011100100100011",  "000011100100111001",  "000011100101001111",  "000011100101100101",  "000011100101111010",  "000011100110010000",  "000011100110100101",  "000011100110111011",  "000011100111010000",  "000011100111100101",  "000011100111111010",  "000011101000001111",  "000011101000100011",  "000011101000111000",  "000011101001001101",  "000011101001100001",  "000011101001110101",  "000011101010001001",  "000011101010011101",  "000011101010110001",  "000011101011000101",  "000011101011011000",  "000011101011101100",  "000011101011111111",  "000011101100010010",  "000011101100100101",  "000011101100111000",  "000011101101001011",  "000011101101011110",  "000011101101110000",  "000011101110000011",  "000011101110010101",  "000011101110100111",  "000011101110111001",  "000011101111001011",  "000011101111011101",  "000011101111101111",  "000011110000000000",  "000011110000010010",  "000011110000100011",  "000011110000110100",  "000011110001000101",  "000011110001010110",  "000011110001100111",  "000011110001110111",  "000011110010001000",  "000011110010011000",  "000011110010101000",  "000011110010111000",  "000011110011001000",  "000011110011011000",  "000011110011101000",  "000011110011110111",  "000011110100000111",  "000011110100010110",  "000011110100100101",  "000011110100110100",  "000011110101000011",  "000011110101010010",  "000011110101100000",  "000011110101101111",  "000011110101111101",  "000011110110001011",  "000011110110011001",  "000011110110100111",  "000011110110110101",  "000011110111000011",  "000011110111010000",  "000011110111011101",  "000011110111101011",  "000011110111111000",  "000011111000000101",  "000011111000010001",  "000011111000011110",  "000011111000101011",  "000011111000110111",  "000011111001000011",  "000011111001001111",  "000011111001011011",  "000011111001100111",  "000011111001110011",  "000011111001111110",  "000011111010001010",  "000011111010010101",  "000011111010100000",  "000011111010101011",  "000011111010110110",  "000011111011000000",  "000011111011001011",  "000011111011010101",  "000011111011100000",  "000011111011101010",  "000011111011110100",  "000011111011111101",  "000011111100000111",  "000011111100010001",  "000011111100011010",  "000011111100100011",  "000011111100101100",  "000011111100110101",  "000011111100111110",  "000011111101000111",  "000011111101001111",  "000011111101011000",  "000011111101100000",  "000011111101101000",  "000011111101110000",  "000011111101111000",  "000011111101111111",  "000011111110000111",  "000011111110001110",  "000011111110010101",  "000011111110011100",  "000011111110100011",  "000011111110101010",  "000011111110110000",  "000011111110110111",  "000011111110111101",  "000011111111000011",  "000011111111001001",  "000011111111001111",  "000011111111010101",  "000011111111011010",  "000011111111100000",  "000011111111100101",  "000011111111101010",  "000011111111101111",  "000011111111110100",  "000011111111111001",  "000011111111111101",  "000100000000000001",  "000100000000000110",  "000100000000001010",  "000100000000001110",  "000100000000010001",  "000100000000010101",  "000100000000011000",  "000100000000011100",  "000100000000011111",  "000100000000100010",  "000100000000100101",  "000100000000100111",  "000100000000101010",  "000100000000101100",  "000100000000101110",  "000100000000110000",  "000100000000110010",  "000100000000110100",  "000100000000110110",  "000100000000110111",  "000100000000111001",  "000100000000111010",  "000100000000111011",  "000100000000111011",  "000100000000111100",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111100",  "000100000000111011",  "000100000000111010",  "000100000000111001",  "000100000000111000",  "000100000000110111",  "000100000000110101",  "000100000000110100",  "000100000000110010",  "000100000000110000",  "000100000000101110",  "000100000000101100",  "000100000000101001",  "000100000000100111",  "000100000000100100",  "000100000000100001",  "000100000000011110",  "000100000000011011",  "000100000000010111",  "000100000000010100",  "000100000000010000",  "000100000000001100",  "000100000000001000",  "000100000000000100",  "000100000000000000",  "000011111111111011",  "000011111111110110",  "000011111111110010",  "000011111111101101",  "000011111111101000",  "000011111111100010",  "000011111111011101",  "000011111111010111",  "000011111111010010",  "000011111111001100",  "000011111111000110",  "000011111110111111",  "000011111110111001",  "000011111110110010",  "000011111110101100",  "000011111110100101",  "000011111110011110",  "000011111110010111",  "000011111110001111",  "000011111110001000",  "000011111110000000",  "000011111101111000",  "000011111101110000",  "000011111101101000",  "000011111101100000",  "000011111101010111",  "000011111101001111",  "000011111101000110",  "000011111100111101",  "000011111100110100",  "000011111100101011",  "000011111100100001",  "000011111100011000",  "000011111100001110",  "000011111100000100",  "000011111011111010",  "000011111011110000",  "000011111011100101",  "000011111011011011",  "000011111011010000",  "000011111011000101",  "000011111010111010",  "000011111010101111",  "000011111010100011",  "000011111010011000",  "000011111010001100",  "000011111010000000",  "000011111001110100",  "000011111001101000",  "000011111001011100",  "000011111001001111",  "000011111001000011",  "000011111000110110",  "000011111000101001",  "000011111000011100",  "000011111000001110",  "000011111000000001",  "000011110111110011",  "000011110111100110",  "000011110111011000",  "000011110111001010",  "000011110110111011",  "000011110110101101",  "000011110110011110",  "000011110110010000",  "000011110110000001",  "000011110101110010",  "000011110101100010",  "000011110101010011",  "000011110101000011",  "000011110100110100",  "000011110100100100",  "000011110100010100",  "000011110100000100",  "000011110011110011",  "000011110011100011",  "000011110011010010",  "000011110011000001",  "000011110010110000",  "000011110010011111",  "000011110010001110",  "000011110001111100",  "000011110001101010",  "000011110001011001",  "000011110001000111",  "000011110000110101",  "000011110000100010",  "000011110000010000",  "000011101111111101",  "000011101111101010",  "000011101111010111",  "000011101111000100",  "000011101110110001",  "000011101110011110",  "000011101110001010",  "000011101101110110",  "000011101101100010",  "000011101101001110",  "000011101100111010",  "000011101100100110",  "000011101100010001",  "000011101011111100",  "000011101011101000",  "000011101011010011",  "000011101010111101",  "000011101010101000",  "000011101010010010",  "000011101001111101",  "000011101001100111",  "000011101001010001",  "000011101000111011",  "000011101000100101",  "000011101000001110",  "000011100111110111",  "000011100111100001",  "000011100111001010",  "000011100110110011",  "000011100110011011",  "000011100110000100",  "000011100101101100",  "000011100101010100",  "000011100100111101",  "000011100100100100",  "000011100100001100",  "000011100011110100",  "000011100011011011",  "000011100011000011",  "000011100010101010",  "000011100010010001",  "000011100001111000",  "000011100001011110",  "000011100001000101",  "000011100000101011",  "000011100000010001",  "000011011111110111",  "000011011111011101",  "000011011111000011",  "000011011110101000",  "000011011110001110",  "000011011101110011",  "000011011101011000",  "000011011100111101",  "000011011100100010",  "000011011100000110",  "000011011011101011",  "000011011011001111",  "000011011010110011",  "000011011010010111",  "000011011001111011",  "000011011001011111",  "000011011001000010",  "000011011000100101",  "000011011000001001",  "000011010111101100",  "000011010111001111",  "000011010110110001",  "000011010110010100",  "000011010101110110",  "000011010101011001",  "000011010100111011",  "000011010100011101",  "000011010011111110",  "000011010011100000",  "000011010011000001",  "000011010010100011",  "000011010010000100",  "000011010001100101",  "000011010001000110",  "000011010000100111",  "000011010000000111",  "000011001111100111",  "000011001111001000",  "000011001110101000",  "000011001110001000",  "000011001101101000",  "000011001101000111",  "000011001100100111",  "000011001100000110",  "000011001011100101",  "000011001011000100",  "000011001010100011",  "000011001010000010",  "000011001001100000",  "000011001000111111",  "000011001000011101",  "000011000111111011",  "000011000111011001",  "000011000110110111",  "000011000110010100",  "000011000101110010",  "000011000101001111",  "000011000100101101",  "000011000100001010",  "000011000011100110",  "000011000011000011",  "000011000010100000",  "000011000001111100",  "000011000001011001",  "000011000000110101",  "000011000000010001",  "000010111111101101",  "000010111111001000",  "000010111110100100",  "000010111101111111",  "000010111101011011",  "000010111100110110",  "000010111100010001",  "000010111011101011",  "000010111011000110",  "000010111010100001",  "000010111001111011",  "000010111001010101",  "000010111000101111",  "000010111000001001",  "000010110111100011",  "000010110110111101",  "000010110110010110",  "000010110101110000",  "000010110101001001",  "000010110100100010",  "000010110011111011",  "000010110011010100",  "000010110010101100",  "000010110010000101",  "000010110001011101",  "000010110000110101",  "000010110000001101",  "000010101111100101",  "000010101110111101",  "000010101110010101",  "000010101101101100",  "000010101101000011",  "000010101100011011",  "000010101011110010",  "000010101011001001",  "000010101010011111",  "000010101001110110",  "000010101001001101",  "000010101000100011",  "000010100111111001",  "000010100111001111",  "000010100110100101",  "000010100101111011",  "000010100101010001",  "000010100100100110",  "000010100011111100",  "000010100011010001",  "000010100010100110",  "000010100001111011",  "000010100001010000",  "000010100000100100",  "000010011111111001",  "000010011111001101",  "000010011110100010",  "000010011101110110",  "000010011101001010",  "000010011100011110",  "000010011011110001",  "000010011011000101",  "000010011010011000",  "000010011001101100",  "000010011000111111",  "000010011000010010",  "000010010111100101",  "000010010110111000",  "000010010110001010",  "000010010101011101",  "000010010100101111",  "000010010100000010",  "000010010011010100",  "000010010010100110",  "000010010001111000",  "000010010001001001",  "000010010000011011",  "000010001111101100",  "000010001110111110",  "000010001110001111",  "000010001101100000",  "000010001100110001",  "000010001100000010",  "000010001011010011",  "000010001010100011",  "000010001001110100",  "000010001001000100",  "000010001000010100",  "000010000111100100",  "000010000110110100",  "000010000110000100",  "000010000101010100",  "000010000100100011",  "000010000011110011",  "000010000011000010",  "000010000010010001",  "000010000001100000",  "000010000000101111",  "000001111111111110",  "000001111111001100",  "000001111110011011",  "000001111101101001",  "000001111100111000",  "000001111100000110",  "000001111011010100",  "000001111010100010",  "000001111001110000",  "000001111000111101",  "000001111000001011",  "000001110111011001",  "000001110110100110",  "000001110101110011",  "000001110101000000",  "000001110100001101",  "000001110011011010",  "000001110010100111",  "000001110001110011",  "000001110001000000",  "000001110000001100",  "000001101111011001",  "000001101110100101",  "000001101101110001",  "000001101100111101",  "000001101100001001",  "000001101011010100",  "000001101010100000",  "000001101001101011",  "000001101000110111",  "000001101000000010",  "000001100111001101",  "000001100110011000",  "000001100101100011",  "000001100100101110",  "000001100011111000",  "000001100011000011",  "000001100010001101",  "000001100001011000",  "000001100000100010",  "000001011111101100",  "000001011110110110",  "000001011110000000",  "000001011101001010",  "000001011100010011",  "000001011011011101",  "000001011010100111",  "000001011001110000",  "000001011000111001",  "000001011000000010",  "000001010111001011",  "000001010110010100",  "000001010101011101",  "000001010100100110",  "000001010011101110",  "000001010010110111",  "000001010001111111",  "000001010001001000",  "000001010000010000",  "000001001111011000",  "000001001110100000",  "000001001101101000",  "000001001100110000",  "000001001011110111",  "000001001010111111",  "000001001010000111",  "000001001001001110",  "000001001000010101",  "000001000111011100",  "000001000110100100",  "000001000101101011",  "000001000100110001",  "000001000011111000",  "000001000010111111",  "000001000010000110",  "000001000001001100",  "000001000000010011",  "000000111111011001",  "000000111110011111",  "000000111101100101",  "000000111100101011",  "000000111011110001",  "000000111010110111",  "000000111001111101",  "000000111001000011",  "000000111000001000",  "000000110111001110",  "000000110110010011",  "000000110101011000",  "000000110100011110",  "000000110011100011",  "000000110010101000",  "000000110001101101",  "000000110000110010",  "000000101111110110",  "000000101110111011",  "000000101110000000",  "000000101101000100",  "000000101100001001",  "000000101011001101",  "000000101010010001",  "000000101001010101",  "000000101000011010",  "000000100111011110",  "000000100110100010",  "000000100101100101",  "000000100100101001",  "000000100011101101",  "000000100010110000",  "000000100001110100",  "000000100000110111",  "000000011111111011",  "000000011110111110",  "000000011110000001",  "000000011101000100",  "000000011100000111",  "000000011011001010",  "000000011010001101",  "000000011001010000",  "000000011000010011",  "000000010111010101",  "000000010110011000",  "000000010101011011",  "000000010100011101",  "000000010011011111",  "000000010010100010",  "000000010001100100",  "000000010000100110",  "000000001111101000",  "000000001110101010",  "000000001101101100",  "000000001100101110",  "000000001011110000",  "000000001010110001",  "000000001001110011",  "000000001000110101",  "000000000111110110",  "000000000110111000",  "000000000101111001",  "000000000100111010",  "000000000011111100",  "000000000010111101",  "000000000001111110",  "000000000000111111"),("000000000000000000",  "111111111111000001",  "111111111110000010",  "111111111101000011",  "111111111100000011",  "111111111011000100",  "111111111010000101",  "111111111001000101",  "111111111000000110",  "111111110111000110",  "111111110110000111",  "111111110101000111",  "111111110100000111",  "111111110011000111",  "111111110010000111",  "111111110001001000",  "111111110000001000",  "111111101111001000",  "111111101110001000",  "111111101101000111",  "111111101100000111",  "111111101011000111",  "111111101010000111",  "111111101001000110",  "111111101000000110",  "111111100111000110",  "111111100110000101",  "111111100101000101",  "111111100100000100",  "111111100011000011",  "111111100010000011",  "111111100001000010",  "111111100000000001",  "111111011111000000",  "111111011101111111",  "111111011100111110",  "111111011011111110",  "111111011010111100",  "111111011001111011",  "111111011000111010",  "111111010111111001",  "111111010110111000",  "111111010101110111",  "111111010100110110",  "111111010011110100",  "111111010010110011",  "111111010001110001",  "111111010000110000",  "111111001111101111",  "111111001110101101",  "111111001101101100",  "111111001100101010",  "111111001011101000",  "111111001010100111",  "111111001001100101",  "111111001000100011",  "111111000111100010",  "111111000110100000",  "111111000101011110",  "111111000100011100",  "111111000011011010",  "111111000010011000",  "111111000001010110",  "111111000000010100",  "111110111111010010",  "111110111110010000",  "111110111101001110",  "111110111100001100",  "111110111011001010",  "111110111010001000",  "111110111001000110",  "111110111000000011",  "111110110111000001",  "111110110101111111",  "111110110100111101",  "111110110011111010",  "111110110010111000",  "111110110001110110",  "111110110000110011",  "111110101111110001",  "111110101110101110",  "111110101101101100",  "111110101100101010",  "111110101011100111",  "111110101010100101",  "111110101001100010",  "111110101000100000",  "111110100111011101",  "111110100110011010",  "111110100101011000",  "111110100100010101",  "111110100011010011",  "111110100010010000",  "111110100001001101",  "111110100000001011",  "111110011111001000",  "111110011110000101",  "111110011101000011",  "111110011100000000",  "111110011010111101",  "111110011001111011",  "111110011000111000",  "111110010111110101",  "111110010110110010",  "111110010101110000",  "111110010100101101",  "111110010011101010",  "111110010010100111",  "111110010001100101",  "111110010000100010",  "111110001111011111",  "111110001110011100",  "111110001101011010",  "111110001100010111",  "111110001011010100",  "111110001010010001",  "111110001001001110",  "111110001000001100",  "111110000111001001",  "111110000110000110",  "111110000101000011",  "111110000100000001",  "111110000010111110",  "111110000001111011",  "111110000000111000",  "111101111111110110",  "111101111110110011",  "111101111101110000",  "111101111100101101",  "111101111011101011",  "111101111010101000",  "111101111001100101",  "111101111000100010",  "111101110111100000",  "111101110110011101",  "111101110101011010",  "111101110100011000",  "111101110011010101",  "111101110010010011",  "111101110001010000",  "111101110000001101",  "111101101111001011",  "111101101110001000",  "111101101101000110",  "111101101100000011",  "111101101011000001",  "111101101001111110",  "111101101000111100",  "111101100111111001",  "111101100110110111",  "111101100101110100",  "111101100100110010",  "111101100011110000",  "111101100010101101",  "111101100001101011",  "111101100000101001",  "111101011111100110",  "111101011110100100",  "111101011101100010",  "111101011100100000",  "111101011011011101",  "111101011010011011",  "111101011001011001",  "111101011000010111",  "111101010111010101",  "111101010110010011",  "111101010101010001",  "111101010100001111",  "111101010011001101",  "111101010010001011",  "111101010001001001",  "111101010000000111",  "111101001111000110",  "111101001110000100",  "111101001101000010",  "111101001100000000",  "111101001010111111",  "111101001001111101",  "111101001000111011",  "111101000111111010",  "111101000110111000",  "111101000101110111",  "111101000100110101",  "111101000011110100",  "111101000010110011",  "111101000001110001",  "111101000000110000",  "111100111111101111",  "111100111110101110",  "111100111101101101",  "111100111100101100",  "111100111011101011",  "111100111010101010",  "111100111001101001",  "111100111000101000",  "111100110111100111",  "111100110110100110",  "111100110101100101",  "111100110100100101",  "111100110011100100",  "111100110010100011",  "111100110001100011",  "111100110000100010",  "111100101111100010",  "111100101110100010",  "111100101101100001",  "111100101100100001",  "111100101011100001",  "111100101010100001",  "111100101001100000",  "111100101000100000",  "111100100111100000",  "111100100110100001",  "111100100101100001",  "111100100100100001",  "111100100011100001",  "111100100010100001",  "111100100001100010",  "111100100000100010",  "111100011111100011",  "111100011110100011",  "111100011101100100",  "111100011100100101",  "111100011011100101",  "111100011010100110",  "111100011001100111",  "111100011000101000",  "111100010111101001",  "111100010110101010",  "111100010101101100",  "111100010100101101",  "111100010011101110",  "111100010010101111",  "111100010001110001",  "111100010000110010",  "111100001111110100",  "111100001110110110",  "111100001101111000",  "111100001100111001",  "111100001011111011",  "111100001010111101",  "111100001001111111",  "111100001001000010",  "111100001000000100",  "111100000111000110",  "111100000110001000",  "111100000101001011",  "111100000100001110",  "111100000011010000",  "111100000010010011",  "111100000001010110",  "111100000000011001",  "111011111111011100",  "111011111110011111",  "111011111101100010",  "111011111100100101",  "111011111011101000",  "111011111010101100",  "111011111001101111",  "111011111000110011",  "111011110111110110",  "111011110110111010",  "111011110101111110",  "111011110101000010",  "111011110100000110",  "111011110011001010",  "111011110010001110",  "111011110001010011",  "111011110000010111",  "111011101111011100",  "111011101110100000",  "111011101101100101",  "111011101100101010",  "111011101011101111",  "111011101010110100",  "111011101001111001",  "111011101000111110",  "111011101000000011",  "111011100111001001",  "111011100110001110",  "111011100101010100",  "111011100100011001",  "111011100011011111",  "111011100010100101",  "111011100001101011",  "111011100000110001",  "111011011111111000",  "111011011110111110",  "111011011110000100",  "111011011101001011",  "111011011100010010",  "111011011011011000",  "111011011010011111",  "111011011001100110",  "111011011000101101",  "111011010111110101",  "111011010110111100",  "111011010110000011",  "111011010101001011",  "111011010100010011",  "111011010011011010",  "111011010010100010",  "111011010001101010",  "111011010000110010",  "111011001111111011",  "111011001111000011",  "111011001110001100",  "111011001101010100",  "111011001100011101",  "111011001011100110",  "111011001010101111",  "111011001001111000",  "111011001001000001",  "111011001000001010",  "111011000111010100",  "111011000110011101",  "111011000101100111",  "111011000100110001",  "111011000011111011",  "111011000011000101",  "111011000010001111",  "111011000001011010",  "111011000000100100",  "111010111111101111",  "111010111110111001",  "111010111110000100",  "111010111101001111",  "111010111100011010",  "111010111011100110",  "111010111010110001",  "111010111001111101",  "111010111001001000",  "111010111000010100",  "111010110111100000",  "111010110110101100",  "111010110101111000",  "111010110101000101",  "111010110100010001",  "111010110011011110",  "111010110010101011",  "111010110001111000",  "111010110001000101",  "111010110000010010",  "111010101111011111",  "111010101110101101",  "111010101101111010",  "111010101101001000",  "111010101100010110",  "111010101011100100",  "111010101010110010",  "111010101010000000",  "111010101001001111",  "111010101000011110",  "111010100111101100",  "111010100110111011",  "111010100110001010",  "111010100101011010",  "111010100100101001",  "111010100011111001",  "111010100011001000",  "111010100010011000",  "111010100001101000",  "111010100000111000",  "111010100000001001",  "111010011111011001",  "111010011110101010",  "111010011101111010",  "111010011101001011",  "111010011100011100",  "111010011011101110",  "111010011010111111",  "111010011010010001",  "111010011001100010",  "111010011000110100",  "111010011000000110",  "111010010111011000",  "111010010110101011",  "111010010101111101",  "111010010101010000",  "111010010100100011",  "111010010011110110",  "111010010011001001",  "111010010010011100",  "111010010001110000",  "111010010001000100",  "111010010000010111",  "111010001111101011",  "111010001111000000",  "111010001110010100",  "111010001101101000",  "111010001100111101",  "111010001100010010",  "111010001011100111",  "111010001010111100",  "111010001010010010",  "111010001001100111",  "111010001000111101",  "111010001000010011",  "111010000111101001",  "111010000110111111",  "111010000110010110",  "111010000101101100",  "111010000101000011",  "111010000100011010",  "111010000011110001",  "111010000011001000",  "111010000010100000",  "111010000001110111",  "111010000001001111",  "111010000000100111",  "111010000000000000",  "111001111111011000",  "111001111110110001",  "111001111110001001",  "111001111101100010",  "111001111100111011",  "111001111100010101",  "111001111011101110",  "111001111011001000",  "111001111010100010",  "111001111001111100",  "111001111001010110",  "111001111000110001",  "111001111000001011",  "111001110111100110",  "111001110111000001",  "111001110110011100",  "111001110101111000",  "111001110101010011",  "111001110100101111",  "111001110100001011",  "111001110011100111",  "111001110011000100",  "111001110010100000",  "111001110001111101",  "111001110001011010",  "111001110000110111",  "111001110000010100",  "111001101111110010",  "111001101111010000",  "111001101110101101",  "111001101110001100",  "111001101101101010",  "111001101101001000",  "111001101100100111",  "111001101100000110",  "111001101011100101",  "111001101011000101",  "111001101010100100",  "111001101010000100",  "111001101001100100",  "111001101001000100",  "111001101000100100",  "111001101000000101",  "111001100111100110",  "111001100111000111",  "111001100110101000",  "111001100110001001",  "111001100101101011",  "111001100101001101",  "111001100100101111",  "111001100100010001",  "111001100011110011",  "111001100011010110",  "111001100010111001",  "111001100010011100",  "111001100001111111",  "111001100001100011",  "111001100001000111",  "111001100000101011",  "111001100000001111",  "111001011111110011",  "111001011111011000",  "111001011110111100",  "111001011110100001",  "111001011110000111",  "111001011101101100",  "111001011101010010",  "111001011100111000",  "111001011100011110",  "111001011100000100",  "111001011011101011",  "111001011011010001",  "111001011010111000",  "111001011010100000",  "111001011010000111",  "111001011001101111",  "111001011001010111",  "111001011000111111",  "111001011000100111",  "111001011000010000",  "111001010111111000",  "111001010111100001",  "111001010111001011",  "111001010110110100",  "111001010110011110",  "111001010110001000",  "111001010101110010",  "111001010101011100",  "111001010101000111",  "111001010100110001",  "111001010100011101",  "111001010100001000",  "111001010011110011",  "111001010011011111",  "111001010011001011",  "111001010010110111",  "111001010010100100",  "111001010010010000",  "111001010001111101",  "111001010001101011",  "111001010001011000",  "111001010001000110",  "111001010000110011",  "111001010000100001",  "111001010000010000",  "111001001111111110",  "111001001111101101",  "111001001111011100",  "111001001111001011",  "111001001110111011",  "111001001110101011",  "111001001110011011",  "111001001110001011",  "111001001101111100",  "111001001101101100",  "111001001101011101",  "111001001101001110",  "111001001101000000",  "111001001100110010",  "111001001100100011",  "111001001100010110",  "111001001100001000",  "111001001011111011",  "111001001011101110",  "111001001011100001",  "111001001011010100",  "111001001011001000",  "111001001010111100",  "111001001010110000",  "111001001010100100",  "111001001010011001",  "111001001010001110",  "111001001010000011",  "111001001001111001",  "111001001001101110",  "111001001001100100",  "111001001001011010",  "111001001001010001",  "111001001001000111",  "111001001000111110",  "111001001000110101",  "111001001000101101",  "111001001000100100",  "111001001000011100",  "111001001000010101",  "111001001000001101",  "111001001000000110",  "111001000111111111",  "111001000111111000",  "111001000111110001",  "111001000111101011",  "111001000111100101",  "111001000111011111",  "111001000111011010",  "111001000111010100",  "111001000111001111",  "111001000111001011",  "111001000111000110",  "111001000111000010",  "111001000110111110",  "111001000110111010",  "111001000110110111",  "111001000110110100",  "111001000110110001",  "111001000110101110",  "111001000110101100",  "111001000110101010",  "111001000110101000",  "111001000110100110",  "111001000110100101",  "111001000110100100",  "111001000110100011",  "111001000110100010",  "111001000110100010",  "111001000110100010",  "111001000110100010",  "111001000110100011",  "111001000110100100",  "111001000110100101",  "111001000110100110",  "111001000110101000",  "111001000110101010",  "111001000110101100",  "111001000110101110",  "111001000110110001",  "111001000110110100",  "111001000110110111",  "111001000110111011",  "111001000110111110",  "111001000111000010",  "111001000111000111",  "111001000111001011",  "111001000111010000",  "111001000111010101",  "111001000111011011",  "111001000111100000",  "111001000111100110",  "111001000111101101",  "111001000111110011",  "111001000111111010",  "111001001000000001",  "111001001000001000",  "111001001000010000",  "111001001000011000",  "111001001000100000",  "111001001000101000",  "111001001000110001",  "111001001000111010",  "111001001001000011",  "111001001001001101",  "111001001001010111",  "111001001001100001",  "111001001001101011",  "111001001001110110",  "111001001010000001",  "111001001010001100",  "111001001010010111",  "111001001010100011",  "111001001010101111",  "111001001010111100",  "111001001011001000",  "111001001011010101",  "111001001011100010",  "111001001011110000",  "111001001011111110",  "111001001100001100",  "111001001100011010",  "111001001100101001",  "111001001100110111",  "111001001101000111",  "111001001101010110",  "111001001101100110",  "111001001101110110",  "111001001110000110",  "111001001110010111",  "111001001110101000",  "111001001110111001",  "111001001111001010",  "111001001111011100",  "111001001111101110",  "111001010000000000",  "111001010000010011",  "111001010000100110",  "111001010000111001",  "111001010001001101",  "111001010001100000",  "111001010001110100",  "111001010010001001",  "111001010010011101",  "111001010010110010",  "111001010011001000",  "111001010011011101",  "111001010011110011",  "111001010100001001",  "111001010100011111",  "111001010100110110",  "111001010101001101",  "111001010101100100",  "111001010101111100",  "111001010110010100",  "111001010110101100",  "111001010111000100",  "111001010111011101",  "111001010111110110",  "111001011000001111",  "111001011000101001",  "111001011001000011",  "111001011001011101",  "111001011001110111",  "111001011010010010",  "111001011010101101",  "111001011011001000",  "111001011011100100",  "111001011100000000",  "111001011100011100",  "111001011100111001",  "111001011101010110",  "111001011101110011",  "111001011110010000",  "111001011110101110",  "111001011111001100",  "111001011111101010",  "111001100000001001",  "111001100000101000",  "111001100001000111",  "111001100001100110",  "111001100010000110",  "111001100010100110",  "111001100011000111",  "111001100011100111",  "111001100100001000",  "111001100100101010",  "111001100101001011",  "111001100101101101",  "111001100110001111",  "111001100110110010",  "111001100111010101",  "111001100111111000",  "111001101000011011",  "111001101000111111",  "111001101001100011",  "111001101010000111",  "111001101010101100",  "111001101011010000",  "111001101011110110",  "111001101100011011",  "111001101101000001",  "111001101101100111",  "111001101110001101",  "111001101110110100",  "111001101111011011",  "111001110000000010",  "111001110000101010",  "111001110001010010",  "111001110001111010",  "111001110010100011",  "111001110011001011",  "111001110011110100",  "111001110100011110",  "111001110101001000",  "111001110101110010",  "111001110110011100",  "111001110111000111",  "111001110111110001",  "111001111000011101",  "111001111001001000",  "111001111001110100",  "111001111010100000",  "111001111011001101",  "111001111011111001",  "111001111100100110",  "111001111101010100",  "111001111110000001",  "111001111110101111",  "111001111111011110",  "111010000000001100",  "111010000000111011",  "111010000001101010",  "111010000010011010",  "111010000011001010",  "111010000011111010",  "111010000100101010",  "111010000101011011",  "111010000110001100",  "111010000110111101",  "111010000111101111",  "111010001000100001",  "111010001001010011",  "111010001010000101",  "111010001010111000",  "111010001011101011",  "111010001100011111",  "111010001101010011",  "111010001110000111",  "111010001110111011",  "111010001111110000",  "111010010000100101",  "111010010001011010",  "111010010010001111",  "111010010011000101",  "111010010011111100",  "111010010100110010",  "111010010101101001",  "111010010110100000",  "111010010111010111",  "111010011000001111",  "111010011001000111",  "111010011010000000",  "111010011010111000",  "111010011011110001",  "111010011100101010",  "111010011101100100",  "111010011110011110",  "111010011111011000",  "111010100000010010",  "111010100001001101",  "111010100010001000",  "111010100011000100",  "111010100011111111",  "111010100100111011",  "111010100101111000",  "111010100110110100",  "111010100111110001",  "111010101000101111",  "111010101001101100",  "111010101010101010",  "111010101011101000",  "111010101100100111",  "111010101101100101",  "111010101110100100",  "111010101111100100",  "111010110000100100",  "111010110001100100",  "111010110010100100",  "111010110011100100",  "111010110100100101",  "111010110101100111",  "111010110110101000",  "111010110111101010",  "111010111000101100",  "111010111001101111",  "111010111010110001",  "111010111011110100",  "111010111100111000",  "111010111101111011",  "111010111110111111",  "111011000000000100",  "111011000001001000",  "111011000010001101",  "111011000011010010",  "111011000100011000",  "111011000101011110",  "111011000110100100",  "111011000111101010",  "111011001000110001",  "111011001001111000",  "111011001010111111",  "111011001100000111",  "111011001101001111",  "111011001110010111",  "111011001111100000",  "111011010000101001",  "111011010001110010",  "111011010010111011",  "111011010100000101",  "111011010101001111",  "111011010110011001",  "111011010111100100",  "111011011000101111",  "111011011001111010",  "111011011011000110",  "111011011100010010",  "111011011101011110",  "111011011110101011",  "111011011111110111",  "111011100001000100",  "111011100010010010",  "111011100011100000",  "111011100100101110",  "111011100101111100",  "111011100111001011",  "111011101000011001",  "111011101001101001",  "111011101010111000",  "111011101100001000",  "111011101101011000",  "111011101110101001",  "111011101111111001",  "111011110001001010",  "111011110010011100",  "111011110011101101",  "111011110100111111",  "111011110110010010",  "111011110111100100",  "111011111000110111",  "111011111010001010",  "111011111011011110",  "111011111100110001",  "111011111110000101",  "111011111111011010",  "111100000000101110",  "111100000010000011",  "111100000011011001",  "111100000100101110",  "111100000110000100",  "111100000111011010",  "111100001000110001",  "111100001010000111",  "111100001011011110",  "111100001100110110",  "111100001110001101",  "111100001111100101",  "111100010000111110",  "111100010010010110",  "111100010011101111",  "111100010101001000",  "111100010110100010",  "111100010111111011",  "111100011001010101",  "111100011010110000",  "111100011100001010",  "111100011101100101",  "111100011111000000",  "111100100000011100",  "111100100001111000",  "111100100011010100",  "111100100100110000",  "111100100110001101",  "111100100111101010",  "111100101001000111",  "111100101010100101",  "111100101100000010",  "111100101101100001",  "111100101110111111",  "111100110000011110",  "111100110001111101",  "111100110011011100",  "111100110100111100",  "111100110110011100",  "111100110111111100",  "111100111001011100",  "111100111010111101",  "111100111100011110",  "111100111101111111",  "111100111111100001",  "111101000001000011",  "111101000010100101",  "111101000100001000",  "111101000101101011",  "111101000111001110",  "111101001000110001",  "111101001010010101",  "111101001011111001",  "111101001101011101",  "111101001111000010",  "111101010000100110",  "111101010010001100",  "111101010011110001",  "111101010101010111",  "111101010110111101",  "111101011000100011",  "111101011010001001",  "111101011011110000",  "111101011101010111",  "111101011110111111",  "111101100000100111",  "111101100010001111",  "111101100011110111",  "111101100101011111",  "111101100111001000",  "111101101000110001",  "111101101010011011",  "111101101100000100",  "111101101101101110",  "111101101111011001",  "111101110001000011",  "111101110010101110",  "111101110100011001",  "111101110110000100",  "111101110111110000",  "111101111001011100",  "111101111011001000",  "111101111100110101",  "111101111110100001",  "111110000000001111",  "111110000001111100",  "111110000011101001",  "111110000101010111",  "111110000111000110",  "111110001000110100",  "111110001010100011",  "111110001100010010",  "111110001110000001",  "111110001111110001",  "111110010001100000",  "111110010011010000",  "111110010101000001",  "111110010110110001",  "111110011000100010",  "111110011010010100",  "111110011100000101",  "111110011101110111",  "111110011111101001",  "111110100001011011",  "111110100011001110",  "111110100101000000",  "111110100110110100",  "111110101000100111",  "111110101010011011",  "111110101100001111",  "111110101110000011",  "111110101111110111",  "111110110001101100",  "111110110011100001",  "111110110101010110",  "111110110111001100",  "111110111001000001",  "111110111010111000",  "111110111100101110",  "111110111110100100",  "111111000000011011",  "111111000010010010",  "111111000100001010",  "111111000110000001",  "111111000111111001",  "111111001001110010",  "111111001011101010",  "111111001101100011",  "111111001111011100",  "111111010001010101",  "111111010011001110",  "111111010101001000",  "111111010111000010",  "111111011000111100",  "111111011010110111",  "111111011100110010",  "111111011110101101",  "111111100000101000",  "111111100010100100",  "111111100100100000",  "111111100110011100",  "111111101000011000",  "111111101010010101",  "111111101100010001",  "111111101110001111",  "111111110000001100",  "111111110010001010",  "111111110100000111",  "111111110110000110",  "111111111000000100",  "111111111010000011",  "111111111100000001",  "111111111110000001"),("000000000000000000",  "000000000010000000",  "000000000100000000",  "000000000110000000",  "000000001000000000",  "000000001010000001",  "000000001100000010",  "000000001110000011",  "000000010000000100",  "000000010010000110",  "000000010100001000",  "000000010110001010",  "000000011000001100",  "000000011010001111",  "000000011100010010",  "000000011110010101",  "000000100000011000",  "000000100010011100",  "000000100100011111",  "000000100110100100",  "000000101000101000",  "000000101010101100",  "000000101100110001",  "000000101110110110",  "000000110000111100",  "000000110011000001",  "000000110101000111",  "000000110111001101",  "000000111001010011",  "000000111011011010",  "000000111101100000",  "000000111111100111",  "000001000001101110",  "000001000011110110",  "000001000101111101",  "000001001000000101",  "000001001010001101",  "000001001100010110",  "000001001110011110",  "000001010000100111",  "000001010010110000",  "000001010100111010",  "000001010111000011",  "000001011001001101",  "000001011011010111",  "000001011101100001",  "000001011111101011",  "000001100001110110",  "000001100100000001",  "000001100110001100",  "000001101000010111",  "000001101010100011",  "000001101100101111",  "000001101110111011",  "000001110001000111",  "000001110011010011",  "000001110101100000",  "000001110111101101",  "000001111001111010",  "000001111100000111",  "000001111110010101",  "000010000000100011",  "000010000010110001",  "000010000100111111",  "000010000111001101",  "000010001001011100",  "000010001011101011",  "000010001101111010",  "000010010000001001",  "000010010010011001",  "000010010100101000",  "000010010110111000",  "000010011001001000",  "000010011011011001",  "000010011101101001",  "000010011111111010",  "000010100010001011",  "000010100100011100",  "000010100110101110",  "000010101000111111",  "000010101011010001",  "000010101101100011",  "000010101111110110",  "000010110010001000",  "000010110100011011",  "000010110110101110",  "000010111001000001",  "000010111011010100",  "000010111101100111",  "000010111111111011",  "000011000010001111",  "000011000100100011",  "000011000110110111",  "000011001001001100",  "000011001011100001",  "000011001101110101",  "000011010000001011",  "000011010010100000",  "000011010100110101",  "000011010111001011",  "000011011001100001",  "000011011011110111",  "000011011110001101",  "000011100000100100",  "000011100010111010",  "000011100101010001",  "000011100111101000",  "000011101001111111",  "000011101100010111",  "000011101110101110",  "000011110001000110",  "000011110011011110",  "000011110101110110",  "000011111000001111",  "000011111010100111",  "000011111101000000",  "000011111111011001",  "000100000001110010",  "000100000100001011",  "000100000110100101",  "000100001000111110",  "000100001011011000",  "000100001101110010",  "000100010000001101",  "000100010010100111",  "000100010101000001",  "000100010111011100",  "000100011001110111",  "000100011100010010",  "000100011110101110",  "000100100001001001",  "000100100011100101",  "000100100110000000",  "000100101000011100",  "000100101010111000",  "000100101101010101",  "000100101111110001",  "000100110010001110",  "000100110100101011",  "000100110111001000",  "000100111001100101",  "000100111100000010",  "000100111110100000",  "000101000000111101",  "000101000011011011",  "000101000101111001",  "000101001000011000",  "000101001010110110",  "000101001101010100",  "000101001111110011",  "000101010010010010",  "000101010100110001",  "000101010111010000",  "000101011001101111",  "000101011100001111",  "000101011110101110",  "000101100001001110",  "000101100011101110",  "000101100110001110",  "000101101000101110",  "000101101011001111",  "000101101101101111",  "000101110000010000",  "000101110010110001",  "000101110101010010",  "000101110111110011",  "000101111010010100",  "000101111100110110",  "000101111111011000",  "000110000001111001",  "000110000100011011",  "000110000110111101",  "000110001001011111",  "000110001100000010",  "000110001110100100",  "000110010001000111",  "000110010011101010",  "000110010110001101",  "000110011000110000",  "000110011011010011",  "000110011101110110",  "000110100000011010",  "000110100010111101",  "000110100101100001",  "000110101000000101",  "000110101010101001",  "000110101101001101",  "000110101111110010",  "000110110010010110",  "000110110100111011",  "000110110111011111",  "000110111010000100",  "000110111100101001",  "000110111111001110",  "000111000001110011",  "000111000100011001",  "000111000110111110",  "000111001001100100",  "000111001100001010",  "000111001110110000",  "000111010001010110",  "000111010011111100",  "000111010110100010",  "000111011001001000",  "000111011011101111",  "000111011110010101",  "000111100000111100",  "000111100011100011",  "000111100110001010",  "000111101000110001",  "000111101011011000",  "000111101101111111",  "000111110000100111",  "000111110011001110",  "000111110101110110",  "000111111000011110",  "000111111011000110",  "000111111101101110",  "001000000000010110",  "001000000010111110",  "001000000101100110",  "001000001000001111",  "001000001010110111",  "001000001101100000",  "001000010000001001",  "001000010010110010",  "001000010101011011",  "001000011000000100",  "001000011010101101",  "001000011101010110",  "001000011111111111",  "001000100010101001",  "001000100101010010",  "001000100111111100",  "001000101010100110",  "001000101101010000",  "001000101111111010",  "001000110010100100",  "001000110101001110",  "001000110111111000",  "001000111010100010",  "001000111101001101",  "001000111111110111",  "001001000010100010",  "001001000101001101",  "001001000111111000",  "001001001010100010",  "001001001101001101",  "001001001111111000",  "001001010010100100",  "001001010101001111",  "001001010111111010",  "001001011010100101",  "001001011101010001",  "001001011111111100",  "001001100010101000",  "001001100101010100",  "001001101000000000",  "001001101010101011",  "001001101101010111",  "001001110000000011",  "001001110010110000",  "001001110101011100",  "001001111000001000",  "001001111010110100",  "001001111101100001",  "001010000000001101",  "001010000010111010",  "001010000101100110",  "001010001000010011",  "001010001011000000",  "001010001101101100",  "001010010000011001",  "001010010011000110",  "001010010101110011",  "001010011000100000",  "001010011011001101",  "001010011101111011",  "001010100000101000",  "001010100011010101",  "001010100110000011",  "001010101000110000",  "001010101011011110",  "001010101110001011",  "001010110000111001",  "001010110011100110",  "001010110110010100",  "001010111001000010",  "001010111011110000",  "001010111110011101",  "001011000001001011",  "001011000011111001",  "001011000110100111",  "001011001001010101",  "001011001100000100",  "001011001110110010",  "001011010001100000",  "001011010100001110",  "001011010110111100",  "001011011001101011",  "001011011100011001",  "001011011111001000",  "001011100001110110",  "001011100100100101",  "001011100111010011",  "001011101010000010",  "001011101100110000",  "001011101111011111",  "001011110010001110",  "001011110100111100",  "001011110111101011",  "001011111010011010",  "001011111101001001",  "001011111111111000",  "001100000010100110",  "001100000101010101",  "001100001000000100",  "001100001010110011",  "001100001101100010",  "001100010000010001",  "001100010011000000",  "001100010101101111",  "001100011000011110",  "001100011011001110",  "001100011101111101",  "001100100000101100",  "001100100011011011",  "001100100110001010",  "001100101000111001",  "001100101011101001",  "001100101110011000",  "001100110001000111",  "001100110011110110",  "001100110110100110",  "001100111001010101",  "001100111100000100",  "001100111110110100",  "001101000001100011",  "001101000100010010",  "001101000111000010",  "001101001001110001",  "001101001100100000",  "001101001111010000",  "001101010001111111",  "001101010100101110",  "001101010111011110",  "001101011010001101",  "001101011100111101",  "001101011111101100",  "001101100010011011",  "001101100101001011",  "001101100111111010",  "001101101010101001",  "001101101101011001",  "001101110000001000",  "001101110010111000",  "001101110101100111",  "001101111000010110",  "001101111011000110",  "001101111101110101",  "001110000000100100",  "001110000011010011",  "001110000110000011",  "001110001000110010",  "001110001011100001",  "001110001110010001",  "001110010001000000",  "001110010011101111",  "001110010110011110",  "001110011001001101",  "001110011011111100",  "001110011110101100",  "001110100001011011",  "001110100100001010",  "001110100110111001",  "001110101001101000",  "001110101100010111",  "001110101111000110",  "001110110001110101",  "001110110100100100",  "001110110111010011",  "001110111010000010",  "001110111100110000",  "001110111111011111",  "001111000010001110",  "001111000100111101",  "001111000111101011",  "001111001010011010",  "001111001101001001",  "001111001111110111",  "001111010010100110",  "001111010101010100",  "001111011000000011",  "001111011010110001",  "001111011101100000",  "001111100000001110",  "001111100010111101",  "001111100101101011",  "001111101000011001",  "001111101011000111",  "001111101101110101",  "001111110000100011",  "001111110011010001",  "001111110101111111",  "001111111000101101",  "001111111011011011",  "001111111110001001",  "010000000000110111",  "010000000011100101",  "010000000110010010",  "010000001001000000",  "010000001011101110",  "010000001110011011",  "010000010001001001",  "010000010011110110",  "010000010110100011",  "010000011001010001",  "010000011011111110",  "010000011110101011",  "010000100001011000",  "010000100100000101",  "010000100110110010",  "010000101001011111",  "010000101100001100",  "010000101110111000",  "010000110001100101",  "010000110100010010",  "010000110110111110",  "010000111001101011",  "010000111100010111",  "010000111111000011",  "010001000001110000",  "010001000100011100",  "010001000111001000",  "010001001001110100",  "010001001100100000",  "010001001111001100",  "010001010001110111",  "010001010100100011",  "010001010111001111",  "010001011001111010",  "010001011100100110",  "010001011111010001",  "010001100001111100",  "010001100100101000",  "010001100111010011",  "010001101001111110",  "010001101100101001",  "010001101111010011",  "010001110001111110",  "010001110100101001",  "010001110111010011",  "010001111001111110",  "010001111100101000",  "010001111111010010",  "010010000001111101",  "010010000100100111",  "010010000111010001",  "010010001001111011",  "010010001100100100",  "010010001111001110",  "010010010001111000",  "010010010100100001",  "010010010111001010",  "010010011001110100",  "010010011100011101",  "010010011111000110",  "010010100001101111",  "010010100100011000",  "010010100111000000",  "010010101001101001",  "010010101100010010",  "010010101110111010",  "010010110001100010",  "010010110100001010",  "010010110110110011",  "010010111001011010",  "010010111100000010",  "010010111110101010",  "010011000001010010",  "010011000011111001",  "010011000110100000",  "010011001001001000",  "010011001011101111",  "010011001110010110",  "010011010000111101",  "010011010011100011",  "010011010110001010",  "010011011000110000",  "010011011011010111",  "010011011101111101",  "010011100000100011",  "010011100011001001",  "010011100101101111",  "010011101000010101",  "010011101010111010",  "010011101101100000",  "010011110000000101",  "010011110010101010",  "010011110101001111",  "010011110111110100",  "010011111010011001",  "010011111100111110",  "010011111111100010",  "010100000010000110",  "010100000100101011",  "010100000111001111",  "010100001001110011",  "010100001100010110",  "010100001110111010",  "010100010001011110",  "010100010100000001",  "010100010110100100",  "010100011001000111",  "010100011011101010",  "010100011110001101",  "010100100000101111",  "010100100011010010",  "010100100101110100",  "010100101000010110",  "010100101010111000",  "010100101101011010",  "010100101111111100",  "010100110010011101",  "010100110100111111",  "010100110111100000",  "010100111010000001",  "010100111100100010",  "010100111111000011",  "010101000001100011",  "010101000100000100",  "010101000110100100",  "010101001001000100",  "010101001011100100",  "010101001110000100",  "010101010000100011",  "010101010011000011",  "010101010101100010",  "010101011000000001",  "010101011010100000",  "010101011100111111",  "010101011111011101",  "010101100001111011",  "010101100100011010",  "010101100110111000",  "010101101001010110",  "010101101011110011",  "010101101110010001",  "010101110000101110",  "010101110011001011",  "010101110101101000",  "010101111000000101",  "010101111010100010",  "010101111100111110",  "010101111111011010",  "010110000001110110",  "010110000100010010",  "010110000110101110",  "010110001001001001",  "010110001011100101",  "010110001110000000",  "010110010000011011",  "010110010010110101",  "010110010101010000",  "010110010111101010",  "010110011010000101",  "010110011100011111",  "010110011110111000",  "010110100001010010",  "010110100011101011",  "010110100110000100",  "010110101000011101",  "010110101010110110",  "010110101101001111",  "010110101111100111",  "010110110001111111",  "010110110100010111",  "010110110110101111",  "010110111001000111",  "010110111011011110",  "010110111101110101",  "010111000000001100",  "010111000010100011",  "010111000100111010",  "010111000111010000",  "010111001001100110",  "010111001011111100",  "010111001110010010",  "010111010000100111",  "010111010010111101",  "010111010101010010",  "010111010111100110",  "010111011001111011",  "010111011100010000",  "010111011110100100",  "010111100000111000",  "010111100011001100",  "010111100101011111",  "010111100111110010",  "010111101010000110",  "010111101100011000",  "010111101110101011",  "010111110000111110",  "010111110011010000",  "010111110101100010",  "010111110111110100",  "010111111010000101",  "010111111100010111",  "010111111110101000",  "011000000000111000",  "011000000011001001",  "011000000101011010",  "011000000111101010",  "011000001001111010",  "011000001100001001",  "011000001110011001",  "011000010000101000",  "011000010010110111",  "011000010101000110",  "011000010111010100",  "011000011001100011",  "011000011011110001",  "011000011101111111",  "011000100000001100",  "011000100010011010",  "011000100100100111",  "011000100110110100",  "011000101001000000",  "011000101011001101",  "011000101101011001",  "011000101111100101",  "011000110001110000",  "011000110011111100",  "011000110110000111",  "011000111000010010",  "011000111010011100",  "011000111100100111",  "011000111110110001",  "011001000000111011",  "011001000011000100",  "011001000101001110",  "011001000111010111",  "011001001001100000",  "011001001011101000",  "011001001101110001",  "011001001111111001",  "011001010010000001",  "011001010100001000",  "011001010110010000",  "011001011000010111",  "011001011010011110",  "011001011100100100",  "011001011110101010",  "011001100000110001",  "011001100010110110",  "011001100100111100",  "011001100111000001",  "011001101001000110",  "011001101011001011",  "011001101101001111",  "011001101111010011",  "011001110001010111",  "011001110011011011",  "011001110101011110",  "011001110111100001",  "011001111001100100",  "011001111011100111",  "011001111101101001",  "011001111111101011",  "011010000001101101",  "011010000011101110",  "011010000101110000",  "011010000111110000",  "011010001001110001",  "011010001011110001",  "011010001101110010",  "011010001111110001",  "011010010001110001",  "011010010011110000",  "011010010101101111",  "011010010111101110",  "011010011001101100",  "011010011011101010",  "011010011101101000",  "011010011111100110",  "011010100001100011",  "011010100011100000",  "011010100101011100",  "011010100111011001",  "011010101001010101",  "011010101011010001",  "011010101101001100",  "011010101111001000",  "011010110001000011",  "011010110010111101",  "011010110100111000",  "011010110110110010",  "011010111000101011",  "011010111010100101",  "011010111100011110",  "011010111110010111",  "011011000000010000",  "011011000010001000",  "011011000100000000",  "011011000101111000",  "011011000111101111",  "011011001001100110",  "011011001011011101",  "011011001101010011",  "011011001111001010",  "011011010000111111",  "011011010010110101",  "011011010100101010",  "011011010110011111",  "011011011000010100",  "011011011010001000",  "011011011011111100",  "011011011101110000",  "011011011111100100",  "011011100001010111",  "011011100011001010",  "011011100100111100",  "011011100110101110",  "011011101000100000",  "011011101010010010",  "011011101100000011",  "011011101101110100",  "011011101111100101",  "011011110001010101",  "011011110011000101",  "011011110100110101",  "011011110110100100",  "011011111000010011",  "011011111010000010",  "011011111011110001",  "011011111101011111",  "011011111111001101",  "011100000000111010",  "011100000010100111",  "011100000100010100",  "011100000110000001",  "011100000111101101",  "011100001001011001",  "011100001011000100",  "011100001100101111",  "011100001110011010",  "011100010000000101",  "011100010001101111",  "011100010011011001",  "011100010101000011",  "011100010110101100",  "011100011000010101",  "011100011001111110",  "011100011011100110",  "011100011101001110",  "011100011110110101",  "011100100000011101",  "011100100010000100",  "011100100011101010",  "011100100101010001",  "011100100110110111",  "011100101000011100",  "011100101010000010",  "011100101011100111",  "011100101101001011",  "011100101110110000",  "011100110000010011",  "011100110001110111",  "011100110011011010",  "011100110100111101",  "011100110110100000",  "011100111000000010",  "011100111001100100",  "011100111011000110",  "011100111100100111",  "011100111110001000",  "011100111111101000",  "011101000001001001",  "011101000010101001",  "011101000100001000",  "011101000101100111",  "011101000111000110",  "011101001000100101",  "011101001010000011",  "011101001011100001",  "011101001100111110",  "011101001110011011",  "011101001111111000",  "011101010001010100",  "011101010010110000",  "011101010100001100",  "011101010101100111",  "011101010111000011",  "011101011000011101",  "011101011001111000",  "011101011011010001",  "011101011100101011",  "011101011110000100",  "011101011111011101",  "011101100000110110",  "011101100010001110",  "011101100011100110",  "011101100100111101",  "011101100110010100",  "011101100111101011",  "011101101001000010",  "011101101010011000",  "011101101011101101",  "011101101101000011",  "011101101110011000",  "011101101111101100",  "011101110001000001",  "011101110010010100",  "011101110011101000",  "011101110100111011",  "011101110110001110",  "011101110111100000",  "011101111000110011",  "011101111010000100",  "011101111011010110",  "011101111100100111",  "011101111101110111",  "011101111111001000",  "011110000000010111",  "011110000001100111",  "011110000010110110",  "011110000100000101",  "011110000101010011",  "011110000110100010",  "011110000111101111",  "011110001000111101",  "011110001010001010",  "011110001011010110",  "011110001100100010",  "011110001101101110",  "011110001110111010",  "011110010000000101",  "011110010001010000",  "011110010010011010",  "011110010011100100",  "011110010100101110",  "011110010101110111",  "011110010111000000",  "011110011000001000",  "011110011001010000",  "011110011010011000",  "011110011011011111",  "011110011100100110",  "011110011101101101",  "011110011110110011",  "011110011111111001",  "011110100000111111",  "011110100010000100",  "011110100011001001",  "011110100100001101",  "011110100101010001",  "011110100110010101",  "011110100111011000",  "011110101000011011",  "011110101001011101",  "011110101010011111",  "011110101011100001",  "011110101100100010",  "011110101101100011",  "011110101110100100",  "011110101111100100",  "011110110000100100",  "011110110001100011",  "011110110010100010",  "011110110011100001",  "011110110100011111",  "011110110101011101",  "011110110110011010",  "011110110111010111",  "011110111000010100",  "011110111001010000",  "011110111010001100",  "011110111011001000",  "011110111100000011",  "011110111100111110",  "011110111101111000",  "011110111110110010",  "011110111111101100",  "011111000000100101",  "011111000001011110",  "011111000010010110",  "011111000011001110",  "011111000100000110",  "011111000100111101",  "011111000101110100",  "011111000110101011",  "011111000111100001",  "011111001000010111",  "011111001001001100",  "011111001010000001",  "011111001010110101",  "011111001011101010",  "011111001100011101",  "011111001101010001",  "011111001110000100",  "011111001110110110",  "011111001111101000",  "011111010000011010",  "011111010001001011",  "011111010001111100",  "011111010010101101",  "011111010011011101",  "011111010100001101",  "011111010100111100",  "011111010101101011",  "011111010110011010",  "011111010111001000",  "011111010111110110",  "011111011000100100",  "011111011001010001",  "011111011001111101",  "011111011010101001",  "011111011011010101",  "011111011100000001",  "011111011100101100",  "011111011101010110",  "011111011110000001",  "011111011110101010",  "011111011111010100",  "011111011111111101",  "011111100000100101",  "011111100001001110",  "011111100001110110",  "011111100010011101",  "011111100011000100",  "011111100011101011",  "011111100100010001",  "011111100100110111",  "011111100101011100",  "011111100110000001",  "011111100110100110",  "011111100111001010",  "011111100111101110",  "011111101000010001",  "011111101000110100",  "011111101001010111",  "011111101001111001",  "011111101010011011",  "011111101010111100",  "011111101011011101",  "011111101011111110",  "011111101100011110",  "011111101100111110",  "011111101101011101",  "011111101101111100",  "011111101110011010",  "011111101110111001",  "011111101111010110",  "011111101111110100",  "011111110000010001",  "011111110000101101",  "011111110001001001",  "011111110001100101",  "011111110010000000",  "011111110010011011",  "011111110010110101",  "011111110011010000",  "011111110011101001",  "011111110100000010",  "011111110100011011",  "011111110100110100",  "011111110101001100",  "011111110101100011",  "011111110101111011",  "011111110110010001",  "011111110110101000",  "011111110110111110",  "011111110111010011",  "011111110111101001",  "011111110111111101",  "011111111000010010",  "011111111000100110",  "011111111000111001",  "011111111001001100",  "011111111001011111",  "011111111001110001",  "011111111010000011",  "011111111010010101",  "011111111010100110",  "011111111010110111",  "011111111011000111",  "011111111011010111",  "011111111011100110",  "011111111011110101",  "011111111100000100",  "011111111100010010",  "011111111100100000",  "011111111100101101",  "011111111100111010",  "011111111101000111",  "011111111101010011",  "011111111101011110",  "011111111101101010",  "011111111101110101",  "011111111101111111",  "011111111110001001",  "011111111110010011",  "011111111110011100",  "011111111110100101",  "011111111110101110",  "011111111110110110",  "011111111110111101",  "011111111111000100",  "011111111111001011",  "011111111111010010",  "011111111111011000",  "011111111111011101",  "011111111111100010",  "011111111111100111",  "011111111111101011",  "011111111111101111",  "011111111111110011",  "011111111111110110",  "011111111111111001",  "011111111111111011",  "011111111111111101",  "011111111111111110",  "011111111111111111",  "011111111111111111"),("011111111111111111",  "011111111111111111",  "011111111111111111",  "011111111111111110",  "011111111111111101",  "011111111111111011",  "011111111111111001",  "011111111111110110",  "011111111111110011",  "011111111111101111",  "011111111111101011",  "011111111111100111",  "011111111111100010",  "011111111111011101",  "011111111111011000",  "011111111111010010",  "011111111111001011",  "011111111111000100",  "011111111110111101",  "011111111110110110",  "011111111110101110",  "011111111110100101",  "011111111110011100",  "011111111110010011",  "011111111110001001",  "011111111101111111",  "011111111101110101",  "011111111101101010",  "011111111101011110",  "011111111101010011",  "011111111101000111",  "011111111100111010",  "011111111100101101",  "011111111100100000",  "011111111100010010",  "011111111100000100",  "011111111011110101",  "011111111011100110",  "011111111011010111",  "011111111011000111",  "011111111010110111",  "011111111010100110",  "011111111010010101",  "011111111010000011",  "011111111001110001",  "011111111001011111",  "011111111001001100",  "011111111000111001",  "011111111000100110",  "011111111000010010",  "011111110111111101",  "011111110111101001",  "011111110111010011",  "011111110110111110",  "011111110110101000",  "011111110110010001",  "011111110101111011",  "011111110101100011",  "011111110101001100",  "011111110100110100",  "011111110100011011",  "011111110100000010",  "011111110011101001",  "011111110011010000",  "011111110010110101",  "011111110010011011",  "011111110010000000",  "011111110001100101",  "011111110001001001",  "011111110000101101",  "011111110000010001",  "011111101111110100",  "011111101111010110",  "011111101110111001",  "011111101110011010",  "011111101101111100",  "011111101101011101",  "011111101100111110",  "011111101100011110",  "011111101011111110",  "011111101011011101",  "011111101010111100",  "011111101010011011",  "011111101001111001",  "011111101001010111",  "011111101000110100",  "011111101000010001",  "011111100111101110",  "011111100111001010",  "011111100110100110",  "011111100110000001",  "011111100101011100",  "011111100100110111",  "011111100100010001",  "011111100011101011",  "011111100011000100",  "011111100010011101",  "011111100001110110",  "011111100001001110",  "011111100000100101",  "011111011111111101",  "011111011111010100",  "011111011110101010",  "011111011110000001",  "011111011101010110",  "011111011100101100",  "011111011100000001",  "011111011011010101",  "011111011010101001",  "011111011001111101",  "011111011001010001",  "011111011000100100",  "011111010111110110",  "011111010111001000",  "011111010110011010",  "011111010101101011",  "011111010100111100",  "011111010100001101",  "011111010011011101",  "011111010010101101",  "011111010001111100",  "011111010001001011",  "011111010000011010",  "011111001111101000",  "011111001110110110",  "011111001110000100",  "011111001101010001",  "011111001100011101",  "011111001011101010",  "011111001010110101",  "011111001010000001",  "011111001001001100",  "011111001000010111",  "011111000111100001",  "011111000110101011",  "011111000101110100",  "011111000100111101",  "011111000100000110",  "011111000011001110",  "011111000010010110",  "011111000001011110",  "011111000000100101",  "011110111111101100",  "011110111110110010",  "011110111101111000",  "011110111100111110",  "011110111100000011",  "011110111011001000",  "011110111010001100",  "011110111001010000",  "011110111000010100",  "011110110111010111",  "011110110110011010",  "011110110101011101",  "011110110100011111",  "011110110011100001",  "011110110010100010",  "011110110001100011",  "011110110000100100",  "011110101111100100",  "011110101110100100",  "011110101101100011",  "011110101100100010",  "011110101011100001",  "011110101010011111",  "011110101001011101",  "011110101000011011",  "011110100111011000",  "011110100110010101",  "011110100101010001",  "011110100100001101",  "011110100011001001",  "011110100010000100",  "011110100000111111",  "011110011111111001",  "011110011110110011",  "011110011101101101",  "011110011100100110",  "011110011011011111",  "011110011010011000",  "011110011001010000",  "011110011000001000",  "011110010111000000",  "011110010101110111",  "011110010100101110",  "011110010011100100",  "011110010010011010",  "011110010001010000",  "011110010000000101",  "011110001110111010",  "011110001101101110",  "011110001100100010",  "011110001011010110",  "011110001010001010",  "011110001000111101",  "011110000111101111",  "011110000110100010",  "011110000101010011",  "011110000100000101",  "011110000010110110",  "011110000001100111",  "011110000000010111",  "011101111111001000",  "011101111101110111",  "011101111100100111",  "011101111011010110",  "011101111010000100",  "011101111000110011",  "011101110111100000",  "011101110110001110",  "011101110100111011",  "011101110011101000",  "011101110010010100",  "011101110001000001",  "011101101111101100",  "011101101110011000",  "011101101101000011",  "011101101011101101",  "011101101010011000",  "011101101001000010",  "011101100111101011",  "011101100110010100",  "011101100100111101",  "011101100011100110",  "011101100010001110",  "011101100000110110",  "011101011111011101",  "011101011110000100",  "011101011100101011",  "011101011011010001",  "011101011001111000",  "011101011000011101",  "011101010111000011",  "011101010101100111",  "011101010100001100",  "011101010010110000",  "011101010001010100",  "011101001111111000",  "011101001110011011",  "011101001100111110",  "011101001011100001",  "011101001010000011",  "011101001000100101",  "011101000111000110",  "011101000101100111",  "011101000100001000",  "011101000010101001",  "011101000001001001",  "011100111111101000",  "011100111110001000",  "011100111100100111",  "011100111011000110",  "011100111001100100",  "011100111000000010",  "011100110110100000",  "011100110100111101",  "011100110011011010",  "011100110001110111",  "011100110000010011",  "011100101110110000",  "011100101101001011",  "011100101011100111",  "011100101010000010",  "011100101000011100",  "011100100110110111",  "011100100101010001",  "011100100011101010",  "011100100010000100",  "011100100000011101",  "011100011110110101",  "011100011101001110",  "011100011011100110",  "011100011001111110",  "011100011000010101",  "011100010110101100",  "011100010101000011",  "011100010011011001",  "011100010001101111",  "011100010000000101",  "011100001110011010",  "011100001100101111",  "011100001011000100",  "011100001001011001",  "011100000111101101",  "011100000110000001",  "011100000100010100",  "011100000010100111",  "011100000000111010",  "011011111111001101",  "011011111101011111",  "011011111011110001",  "011011111010000010",  "011011111000010011",  "011011110110100100",  "011011110100110101",  "011011110011000101",  "011011110001010101",  "011011101111100101",  "011011101101110100",  "011011101100000011",  "011011101010010010",  "011011101000100000",  "011011100110101110",  "011011100100111100",  "011011100011001010",  "011011100001010111",  "011011011111100100",  "011011011101110000",  "011011011011111100",  "011011011010001000",  "011011011000010100",  "011011010110011111",  "011011010100101010",  "011011010010110101",  "011011010000111111",  "011011001111001010",  "011011001101010011",  "011011001011011101",  "011011001001100110",  "011011000111101111",  "011011000101111000",  "011011000100000000",  "011011000010001000",  "011011000000010000",  "011010111110010111",  "011010111100011110",  "011010111010100101",  "011010111000101011",  "011010110110110010",  "011010110100111000",  "011010110010111101",  "011010110001000011",  "011010101111001000",  "011010101101001100",  "011010101011010001",  "011010101001010101",  "011010100111011001",  "011010100101011100",  "011010100011100000",  "011010100001100011",  "011010011111100110",  "011010011101101000",  "011010011011101010",  "011010011001101100",  "011010010111101110",  "011010010101101111",  "011010010011110000",  "011010010001110001",  "011010001111110001",  "011010001101110010",  "011010001011110001",  "011010001001110001",  "011010000111110000",  "011010000101110000",  "011010000011101110",  "011010000001101101",  "011001111111101011",  "011001111101101001",  "011001111011100111",  "011001111001100100",  "011001110111100001",  "011001110101011110",  "011001110011011011",  "011001110001010111",  "011001101111010011",  "011001101101001111",  "011001101011001011",  "011001101001000110",  "011001100111000001",  "011001100100111100",  "011001100010110110",  "011001100000110001",  "011001011110101010",  "011001011100100100",  "011001011010011110",  "011001011000010111",  "011001010110010000",  "011001010100001000",  "011001010010000001",  "011001001111111001",  "011001001101110001",  "011001001011101000",  "011001001001100000",  "011001000111010111",  "011001000101001110",  "011001000011000100",  "011001000000111011",  "011000111110110001",  "011000111100100111",  "011000111010011100",  "011000111000010010",  "011000110110000111",  "011000110011111100",  "011000110001110000",  "011000101111100101",  "011000101101011001",  "011000101011001101",  "011000101001000000",  "011000100110110100",  "011000100100100111",  "011000100010011010",  "011000100000001100",  "011000011101111111",  "011000011011110001",  "011000011001100011",  "011000010111010100",  "011000010101000110",  "011000010010110111",  "011000010000101000",  "011000001110011001",  "011000001100001001",  "011000001001111010",  "011000000111101010",  "011000000101011010",  "011000000011001001",  "011000000000111000",  "010111111110101000",  "010111111100010111",  "010111111010000101",  "010111110111110100",  "010111110101100010",  "010111110011010000",  "010111110000111110",  "010111101110101011",  "010111101100011000",  "010111101010000110",  "010111100111110010",  "010111100101011111",  "010111100011001100",  "010111100000111000",  "010111011110100100",  "010111011100010000",  "010111011001111011",  "010111010111100110",  "010111010101010010",  "010111010010111101",  "010111010000100111",  "010111001110010010",  "010111001011111100",  "010111001001100110",  "010111000111010000",  "010111000100111010",  "010111000010100011",  "010111000000001100",  "010110111101110101",  "010110111011011110",  "010110111001000111",  "010110110110101111",  "010110110100010111",  "010110110001111111",  "010110101111100111",  "010110101101001111",  "010110101010110110",  "010110101000011101",  "010110100110000100",  "010110100011101011",  "010110100001010010",  "010110011110111000",  "010110011100011111",  "010110011010000101",  "010110010111101010",  "010110010101010000",  "010110010010110101",  "010110010000011011",  "010110001110000000",  "010110001011100101",  "010110001001001001",  "010110000110101110",  "010110000100010010",  "010110000001110110",  "010101111111011010",  "010101111100111110",  "010101111010100010",  "010101111000000101",  "010101110101101000",  "010101110011001011",  "010101110000101110",  "010101101110010001",  "010101101011110011",  "010101101001010110",  "010101100110111000",  "010101100100011010",  "010101100001111011",  "010101011111011101",  "010101011100111111",  "010101011010100000",  "010101011000000001",  "010101010101100010",  "010101010011000011",  "010101010000100011",  "010101001110000100",  "010101001011100100",  "010101001001000100",  "010101000110100100",  "010101000100000100",  "010101000001100011",  "010100111111000011",  "010100111100100010",  "010100111010000001",  "010100110111100000",  "010100110100111111",  "010100110010011101",  "010100101111111100",  "010100101101011010",  "010100101010111000",  "010100101000010110",  "010100100101110100",  "010100100011010010",  "010100100000101111",  "010100011110001101",  "010100011011101010",  "010100011001000111",  "010100010110100100",  "010100010100000001",  "010100010001011110",  "010100001110111010",  "010100001100010110",  "010100001001110011",  "010100000111001111",  "010100000100101011",  "010100000010000110",  "010011111111100010",  "010011111100111110",  "010011111010011001",  "010011110111110100",  "010011110101001111",  "010011110010101010",  "010011110000000101",  "010011101101100000",  "010011101010111010",  "010011101000010101",  "010011100101101111",  "010011100011001001",  "010011100000100011",  "010011011101111101",  "010011011011010111",  "010011011000110000",  "010011010110001010",  "010011010011100011",  "010011010000111101",  "010011001110010110",  "010011001011101111",  "010011001001001000",  "010011000110100000",  "010011000011111001",  "010011000001010010",  "010010111110101010",  "010010111100000010",  "010010111001011010",  "010010110110110011",  "010010110100001010",  "010010110001100010",  "010010101110111010",  "010010101100010010",  "010010101001101001",  "010010100111000000",  "010010100100011000",  "010010100001101111",  "010010011111000110",  "010010011100011101",  "010010011001110100",  "010010010111001010",  "010010010100100001",  "010010010001111000",  "010010001111001110",  "010010001100100100",  "010010001001111011",  "010010000111010001",  "010010000100100111",  "010010000001111101",  "010001111111010010",  "010001111100101000",  "010001111001111110",  "010001110111010011",  "010001110100101001",  "010001110001111110",  "010001101111010011",  "010001101100101001",  "010001101001111110",  "010001100111010011",  "010001100100101000",  "010001100001111100",  "010001011111010001",  "010001011100100110",  "010001011001111010",  "010001010111001111",  "010001010100100011",  "010001010001110111",  "010001001111001100",  "010001001100100000",  "010001001001110100",  "010001000111001000",  "010001000100011100",  "010001000001110000",  "010000111111000011",  "010000111100010111",  "010000111001101011",  "010000110110111110",  "010000110100010010",  "010000110001100101",  "010000101110111000",  "010000101100001100",  "010000101001011111",  "010000100110110010",  "010000100100000101",  "010000100001011000",  "010000011110101011",  "010000011011111110",  "010000011001010001",  "010000010110100011",  "010000010011110110",  "010000010001001001",  "010000001110011011",  "010000001011101110",  "010000001001000000",  "010000000110010010",  "010000000011100101",  "010000000000110111",  "001111111110001001",  "001111111011011011",  "001111111000101101",  "001111110101111111",  "001111110011010001",  "001111110000100011",  "001111101101110101",  "001111101011000111",  "001111101000011001",  "001111100101101011",  "001111100010111101",  "001111100000001110",  "001111011101100000",  "001111011010110001",  "001111011000000011",  "001111010101010100",  "001111010010100110",  "001111001111110111",  "001111001101001001",  "001111001010011010",  "001111000111101011",  "001111000100111101",  "001111000010001110",  "001110111111011111",  "001110111100110000",  "001110111010000010",  "001110110111010011",  "001110110100100100",  "001110110001110101",  "001110101111000110",  "001110101100010111",  "001110101001101000",  "001110100110111001",  "001110100100001010",  "001110100001011011",  "001110011110101100",  "001110011011111100",  "001110011001001101",  "001110010110011110",  "001110010011101111",  "001110010001000000",  "001110001110010001",  "001110001011100001",  "001110001000110010",  "001110000110000011",  "001110000011010011",  "001110000000100100",  "001101111101110101",  "001101111011000110",  "001101111000010110",  "001101110101100111",  "001101110010111000",  "001101110000001000",  "001101101101011001",  "001101101010101001",  "001101100111111010",  "001101100101001011",  "001101100010011011",  "001101011111101100",  "001101011100111101",  "001101011010001101",  "001101010111011110",  "001101010100101110",  "001101010001111111",  "001101001111010000",  "001101001100100000",  "001101001001110001",  "001101000111000010",  "001101000100010010",  "001101000001100011",  "001100111110110100",  "001100111100000100",  "001100111001010101",  "001100110110100110",  "001100110011110110",  "001100110001000111",  "001100101110011000",  "001100101011101001",  "001100101000111001",  "001100100110001010",  "001100100011011011",  "001100100000101100",  "001100011101111101",  "001100011011001110",  "001100011000011110",  "001100010101101111",  "001100010011000000",  "001100010000010001",  "001100001101100010",  "001100001010110011",  "001100001000000100",  "001100000101010101",  "001100000010100110",  "001011111111111000",  "001011111101001001",  "001011111010011010",  "001011110111101011",  "001011110100111100",  "001011110010001110",  "001011101111011111",  "001011101100110000",  "001011101010000010",  "001011100111010011",  "001011100100100101",  "001011100001110110",  "001011011111001000",  "001011011100011001",  "001011011001101011",  "001011010110111100",  "001011010100001110",  "001011010001100000",  "001011001110110010",  "001011001100000100",  "001011001001010101",  "001011000110100111",  "001011000011111001",  "001011000001001011",  "001010111110011101",  "001010111011110000",  "001010111001000010",  "001010110110010100",  "001010110011100110",  "001010110000111001",  "001010101110001011",  "001010101011011110",  "001010101000110000",  "001010100110000011",  "001010100011010101",  "001010100000101000",  "001010011101111011",  "001010011011001101",  "001010011000100000",  "001010010101110011",  "001010010011000110",  "001010010000011001",  "001010001101101100",  "001010001011000000",  "001010001000010011",  "001010000101100110",  "001010000010111010",  "001010000000001101",  "001001111101100001",  "001001111010110100",  "001001111000001000",  "001001110101011100",  "001001110010110000",  "001001110000000011",  "001001101101010111",  "001001101010101011",  "001001101000000000",  "001001100101010100",  "001001100010101000",  "001001011111111100",  "001001011101010001",  "001001011010100101",  "001001010111111010",  "001001010101001111",  "001001010010100100",  "001001001111111000",  "001001001101001101",  "001001001010100010",  "001001000111111000",  "001001000101001101",  "001001000010100010",  "001000111111110111",  "001000111101001101",  "001000111010100010",  "001000110111111000",  "001000110101001110",  "001000110010100100",  "001000101111111010",  "001000101101010000",  "001000101010100110",  "001000100111111100",  "001000100101010010",  "001000100010101001",  "001000011111111111",  "001000011101010110",  "001000011010101101",  "001000011000000100",  "001000010101011011",  "001000010010110010",  "001000010000001001",  "001000001101100000",  "001000001010110111",  "001000001000001111",  "001000000101100110",  "001000000010111110",  "001000000000010110",  "000111111101101110",  "000111111011000110",  "000111111000011110",  "000111110101110110",  "000111110011001110",  "000111110000100111",  "000111101101111111",  "000111101011011000",  "000111101000110001",  "000111100110001010",  "000111100011100011",  "000111100000111100",  "000111011110010101",  "000111011011101111",  "000111011001001000",  "000111010110100010",  "000111010011111100",  "000111010001010110",  "000111001110110000",  "000111001100001010",  "000111001001100100",  "000111000110111110",  "000111000100011001",  "000111000001110011",  "000110111111001110",  "000110111100101001",  "000110111010000100",  "000110110111011111",  "000110110100111011",  "000110110010010110",  "000110101111110010",  "000110101101001101",  "000110101010101001",  "000110101000000101",  "000110100101100001",  "000110100010111101",  "000110100000011010",  "000110011101110110",  "000110011011010011",  "000110011000110000",  "000110010110001101",  "000110010011101010",  "000110010001000111",  "000110001110100100",  "000110001100000010",  "000110001001011111",  "000110000110111101",  "000110000100011011",  "000110000001111001",  "000101111111011000",  "000101111100110110",  "000101111010010100",  "000101110111110011",  "000101110101010010",  "000101110010110001",  "000101110000010000",  "000101101101101111",  "000101101011001111",  "000101101000101110",  "000101100110001110",  "000101100011101110",  "000101100001001110",  "000101011110101110",  "000101011100001111",  "000101011001101111",  "000101010111010000",  "000101010100110001",  "000101010010010010",  "000101001111110011",  "000101001101010100",  "000101001010110110",  "000101001000011000",  "000101000101111001",  "000101000011011011",  "000101000000111101",  "000100111110100000",  "000100111100000010",  "000100111001100101",  "000100110111001000",  "000100110100101011",  "000100110010001110",  "000100101111110001",  "000100101101010101",  "000100101010111000",  "000100101000011100",  "000100100110000000",  "000100100011100101",  "000100100001001001",  "000100011110101110",  "000100011100010010",  "000100011001110111",  "000100010111011100",  "000100010101000001",  "000100010010100111",  "000100010000001101",  "000100001101110010",  "000100001011011000",  "000100001000111110",  "000100000110100101",  "000100000100001011",  "000100000001110010",  "000011111111011001",  "000011111101000000",  "000011111010100111",  "000011111000001111",  "000011110101110110",  "000011110011011110",  "000011110001000110",  "000011101110101110",  "000011101100010111",  "000011101001111111",  "000011100111101000",  "000011100101010001",  "000011100010111010",  "000011100000100100",  "000011011110001101",  "000011011011110111",  "000011011001100001",  "000011010111001011",  "000011010100110101",  "000011010010100000",  "000011010000001011",  "000011001101110101",  "000011001011100001",  "000011001001001100",  "000011000110110111",  "000011000100100011",  "000011000010001111",  "000010111111111011",  "000010111101100111",  "000010111011010100",  "000010111001000001",  "000010110110101110",  "000010110100011011",  "000010110010001000",  "000010101111110110",  "000010101101100011",  "000010101011010001",  "000010101000111111",  "000010100110101110",  "000010100100011100",  "000010100010001011",  "000010011111111010",  "000010011101101001",  "000010011011011001",  "000010011001001000",  "000010010110111000",  "000010010100101000",  "000010010010011001",  "000010010000001001",  "000010001101111010",  "000010001011101011",  "000010001001011100",  "000010000111001101",  "000010000100111111",  "000010000010110001",  "000010000000100011",  "000001111110010101",  "000001111100000111",  "000001111001111010",  "000001110111101101",  "000001110101100000",  "000001110011010011",  "000001110001000111",  "000001101110111011",  "000001101100101111",  "000001101010100011",  "000001101000010111",  "000001100110001100",  "000001100100000001",  "000001100001110110",  "000001011111101011",  "000001011101100001",  "000001011011010111",  "000001011001001101",  "000001010111000011",  "000001010100111010",  "000001010010110000",  "000001010000100111",  "000001001110011110",  "000001001100010110",  "000001001010001101",  "000001001000000101",  "000001000101111101",  "000001000011110110",  "000001000001101110",  "000000111111100111",  "000000111101100000",  "000000111011011010",  "000000111001010011",  "000000110111001101",  "000000110101000111",  "000000110011000001",  "000000110000111100",  "000000101110110110",  "000000101100110001",  "000000101010101100",  "000000101000101000",  "000000100110100100",  "000000100100011111",  "000000100010011100",  "000000100000011000",  "000000011110010101",  "000000011100010010",  "000000011010001111",  "000000011000001100",  "000000010110001010",  "000000010100001000",  "000000010010000110",  "000000010000000100",  "000000001110000011",  "000000001100000010",  "000000001010000001",  "000000001000000000",  "000000000110000000",  "000000000100000000",  "000000000010000000"),("000000000000000000",  "111111111110000001",  "111111111100000001",  "111111111010000011",  "111111111000000100",  "111111110110000110",  "111111110100000111",  "111111110010001010",  "111111110000001100",  "111111101110001111",  "111111101100010001",  "111111101010010101",  "111111101000011000",  "111111100110011100",  "111111100100100000",  "111111100010100100",  "111111100000101000",  "111111011110101101",  "111111011100110010",  "111111011010110111",  "111111011000111100",  "111111010111000010",  "111111010101001000",  "111111010011001110",  "111111010001010101",  "111111001111011100",  "111111001101100011",  "111111001011101010",  "111111001001110010",  "111111000111111001",  "111111000110000001",  "111111000100001010",  "111111000010010010",  "111111000000011011",  "111110111110100100",  "111110111100101110",  "111110111010111000",  "111110111001000001",  "111110110111001100",  "111110110101010110",  "111110110011100001",  "111110110001101100",  "111110101111110111",  "111110101110000011",  "111110101100001111",  "111110101010011011",  "111110101000100111",  "111110100110110100",  "111110100101000000",  "111110100011001110",  "111110100001011011",  "111110011111101001",  "111110011101110111",  "111110011100000101",  "111110011010010100",  "111110011000100010",  "111110010110110001",  "111110010101000001",  "111110010011010000",  "111110010001100000",  "111110001111110001",  "111110001110000001",  "111110001100010010",  "111110001010100011",  "111110001000110100",  "111110000111000110",  "111110000101010111",  "111110000011101001",  "111110000001111100",  "111110000000001111",  "111101111110100001",  "111101111100110101",  "111101111011001000",  "111101111001011100",  "111101110111110000",  "111101110110000100",  "111101110100011001",  "111101110010101110",  "111101110001000011",  "111101101111011001",  "111101101101101110",  "111101101100000100",  "111101101010011011",  "111101101000110001",  "111101100111001000",  "111101100101011111",  "111101100011110111",  "111101100010001111",  "111101100000100111",  "111101011110111111",  "111101011101010111",  "111101011011110000",  "111101011010001001",  "111101011000100011",  "111101010110111101",  "111101010101010111",  "111101010011110001",  "111101010010001100",  "111101010000100110",  "111101001111000010",  "111101001101011101",  "111101001011111001",  "111101001010010101",  "111101001000110001",  "111101000111001110",  "111101000101101011",  "111101000100001000",  "111101000010100101",  "111101000001000011",  "111100111111100001",  "111100111101111111",  "111100111100011110",  "111100111010111101",  "111100111001011100",  "111100110111111100",  "111100110110011100",  "111100110100111100",  "111100110011011100",  "111100110001111101",  "111100110000011110",  "111100101110111111",  "111100101101100001",  "111100101100000010",  "111100101010100101",  "111100101001000111",  "111100100111101010",  "111100100110001101",  "111100100100110000",  "111100100011010100",  "111100100001111000",  "111100100000011100",  "111100011111000000",  "111100011101100101",  "111100011100001010",  "111100011010110000",  "111100011001010101",  "111100010111111011",  "111100010110100010",  "111100010101001000",  "111100010011101111",  "111100010010010110",  "111100010000111110",  "111100001111100101",  "111100001110001101",  "111100001100110110",  "111100001011011110",  "111100001010000111",  "111100001000110001",  "111100000111011010",  "111100000110000100",  "111100000100101110",  "111100000011011001",  "111100000010000011",  "111100000000101110",  "111011111111011010",  "111011111110000101",  "111011111100110001",  "111011111011011110",  "111011111010001010",  "111011111000110111",  "111011110111100100",  "111011110110010010",  "111011110100111111",  "111011110011101101",  "111011110010011100",  "111011110001001010",  "111011101111111001",  "111011101110101001",  "111011101101011000",  "111011101100001000",  "111011101010111000",  "111011101001101001",  "111011101000011001",  "111011100111001011",  "111011100101111100",  "111011100100101110",  "111011100011100000",  "111011100010010010",  "111011100001000100",  "111011011111110111",  "111011011110101011",  "111011011101011110",  "111011011100010010",  "111011011011000110",  "111011011001111010",  "111011011000101111",  "111011010111100100",  "111011010110011001",  "111011010101001111",  "111011010100000101",  "111011010010111011",  "111011010001110010",  "111011010000101001",  "111011001111100000",  "111011001110010111",  "111011001101001111",  "111011001100000111",  "111011001010111111",  "111011001001111000",  "111011001000110001",  "111011000111101010",  "111011000110100100",  "111011000101011110",  "111011000100011000",  "111011000011010010",  "111011000010001101",  "111011000001001000",  "111011000000000100",  "111010111110111111",  "111010111101111011",  "111010111100111000",  "111010111011110100",  "111010111010110001",  "111010111001101111",  "111010111000101100",  "111010110111101010",  "111010110110101000",  "111010110101100111",  "111010110100100101",  "111010110011100100",  "111010110010100100",  "111010110001100100",  "111010110000100100",  "111010101111100100",  "111010101110100100",  "111010101101100101",  "111010101100100111",  "111010101011101000",  "111010101010101010",  "111010101001101100",  "111010101000101111",  "111010100111110001",  "111010100110110100",  "111010100101111000",  "111010100100111011",  "111010100011111111",  "111010100011000100",  "111010100010001000",  "111010100001001101",  "111010100000010010",  "111010011111011000",  "111010011110011110",  "111010011101100100",  "111010011100101010",  "111010011011110001",  "111010011010111000",  "111010011010000000",  "111010011001000111",  "111010011000001111",  "111010010111010111",  "111010010110100000",  "111010010101101001",  "111010010100110010",  "111010010011111100",  "111010010011000101",  "111010010010001111",  "111010010001011010",  "111010010000100101",  "111010001111110000",  "111010001110111011",  "111010001110000111",  "111010001101010011",  "111010001100011111",  "111010001011101011",  "111010001010111000",  "111010001010000101",  "111010001001010011",  "111010001000100001",  "111010000111101111",  "111010000110111101",  "111010000110001100",  "111010000101011011",  "111010000100101010",  "111010000011111010",  "111010000011001010",  "111010000010011010",  "111010000001101010",  "111010000000111011",  "111010000000001100",  "111001111111011110",  "111001111110101111",  "111001111110000001",  "111001111101010100",  "111001111100100110",  "111001111011111001",  "111001111011001101",  "111001111010100000",  "111001111001110100",  "111001111001001000",  "111001111000011101",  "111001110111110001",  "111001110111000111",  "111001110110011100",  "111001110101110010",  "111001110101001000",  "111001110100011110",  "111001110011110100",  "111001110011001011",  "111001110010100011",  "111001110001111010",  "111001110001010010",  "111001110000101010",  "111001110000000010",  "111001101111011011",  "111001101110110100",  "111001101110001101",  "111001101101100111",  "111001101101000001",  "111001101100011011",  "111001101011110110",  "111001101011010000",  "111001101010101100",  "111001101010000111",  "111001101001100011",  "111001101000111111",  "111001101000011011",  "111001100111111000",  "111001100111010101",  "111001100110110010",  "111001100110001111",  "111001100101101101",  "111001100101001011",  "111001100100101010",  "111001100100001000",  "111001100011100111",  "111001100011000111",  "111001100010100110",  "111001100010000110",  "111001100001100110",  "111001100001000111",  "111001100000101000",  "111001100000001001",  "111001011111101010",  "111001011111001100",  "111001011110101110",  "111001011110010000",  "111001011101110011",  "111001011101010110",  "111001011100111001",  "111001011100011100",  "111001011100000000",  "111001011011100100",  "111001011011001000",  "111001011010101101",  "111001011010010010",  "111001011001110111",  "111001011001011101",  "111001011001000011",  "111001011000101001",  "111001011000001111",  "111001010111110110",  "111001010111011101",  "111001010111000100",  "111001010110101100",  "111001010110010100",  "111001010101111100",  "111001010101100100",  "111001010101001101",  "111001010100110110",  "111001010100011111",  "111001010100001001",  "111001010011110011",  "111001010011011101",  "111001010011001000",  "111001010010110010",  "111001010010011101",  "111001010010001001",  "111001010001110100",  "111001010001100000",  "111001010001001101",  "111001010000111001",  "111001010000100110",  "111001010000010011",  "111001010000000000",  "111001001111101110",  "111001001111011100",  "111001001111001010",  "111001001110111001",  "111001001110101000",  "111001001110010111",  "111001001110000110",  "111001001101110110",  "111001001101100110",  "111001001101010110",  "111001001101000111",  "111001001100110111",  "111001001100101001",  "111001001100011010",  "111001001100001100",  "111001001011111110",  "111001001011110000",  "111001001011100010",  "111001001011010101",  "111001001011001000",  "111001001010111100",  "111001001010101111",  "111001001010100011",  "111001001010010111",  "111001001010001100",  "111001001010000001",  "111001001001110110",  "111001001001101011",  "111001001001100001",  "111001001001010111",  "111001001001001101",  "111001001001000011",  "111001001000111010",  "111001001000110001",  "111001001000101000",  "111001001000100000",  "111001001000011000",  "111001001000010000",  "111001001000001000",  "111001001000000001",  "111001000111111010",  "111001000111110011",  "111001000111101101",  "111001000111100110",  "111001000111100000",  "111001000111011011",  "111001000111010101",  "111001000111010000",  "111001000111001011",  "111001000111000111",  "111001000111000010",  "111001000110111110",  "111001000110111011",  "111001000110110111",  "111001000110110100",  "111001000110110001",  "111001000110101110",  "111001000110101100",  "111001000110101010",  "111001000110101000",  "111001000110100110",  "111001000110100101",  "111001000110100100",  "111001000110100011",  "111001000110100010",  "111001000110100010",  "111001000110100010",  "111001000110100010",  "111001000110100011",  "111001000110100100",  "111001000110100101",  "111001000110100110",  "111001000110101000",  "111001000110101010",  "111001000110101100",  "111001000110101110",  "111001000110110001",  "111001000110110100",  "111001000110110111",  "111001000110111010",  "111001000110111110",  "111001000111000010",  "111001000111000110",  "111001000111001011",  "111001000111001111",  "111001000111010100",  "111001000111011010",  "111001000111011111",  "111001000111100101",  "111001000111101011",  "111001000111110001",  "111001000111111000",  "111001000111111111",  "111001001000000110",  "111001001000001101",  "111001001000010101",  "111001001000011100",  "111001001000100100",  "111001001000101101",  "111001001000110101",  "111001001000111110",  "111001001001000111",  "111001001001010001",  "111001001001011010",  "111001001001100100",  "111001001001101110",  "111001001001111001",  "111001001010000011",  "111001001010001110",  "111001001010011001",  "111001001010100100",  "111001001010110000",  "111001001010111100",  "111001001011001000",  "111001001011010100",  "111001001011100001",  "111001001011101110",  "111001001011111011",  "111001001100001000",  "111001001100010110",  "111001001100100011",  "111001001100110010",  "111001001101000000",  "111001001101001110",  "111001001101011101",  "111001001101101100",  "111001001101111100",  "111001001110001011",  "111001001110011011",  "111001001110101011",  "111001001110111011",  "111001001111001011",  "111001001111011100",  "111001001111101101",  "111001001111111110",  "111001010000010000",  "111001010000100001",  "111001010000110011",  "111001010001000110",  "111001010001011000",  "111001010001101011",  "111001010001111101",  "111001010010010000",  "111001010010100100",  "111001010010110111",  "111001010011001011",  "111001010011011111",  "111001010011110011",  "111001010100001000",  "111001010100011101",  "111001010100110001",  "111001010101000111",  "111001010101011100",  "111001010101110010",  "111001010110001000",  "111001010110011110",  "111001010110110100",  "111001010111001011",  "111001010111100001",  "111001010111111000",  "111001011000010000",  "111001011000100111",  "111001011000111111",  "111001011001010111",  "111001011001101111",  "111001011010000111",  "111001011010100000",  "111001011010111000",  "111001011011010001",  "111001011011101011",  "111001011100000100",  "111001011100011110",  "111001011100111000",  "111001011101010010",  "111001011101101100",  "111001011110000111",  "111001011110100001",  "111001011110111100",  "111001011111011000",  "111001011111110011",  "111001100000001111",  "111001100000101011",  "111001100001000111",  "111001100001100011",  "111001100001111111",  "111001100010011100",  "111001100010111001",  "111001100011010110",  "111001100011110011",  "111001100100010001",  "111001100100101111",  "111001100101001101",  "111001100101101011",  "111001100110001001",  "111001100110101000",  "111001100111000111",  "111001100111100110",  "111001101000000101",  "111001101000100100",  "111001101001000100",  "111001101001100100",  "111001101010000100",  "111001101010100100",  "111001101011000101",  "111001101011100101",  "111001101100000110",  "111001101100100111",  "111001101101001000",  "111001101101101010",  "111001101110001100",  "111001101110101101",  "111001101111010000",  "111001101111110010",  "111001110000010100",  "111001110000110111",  "111001110001011010",  "111001110001111101",  "111001110010100000",  "111001110011000100",  "111001110011100111",  "111001110100001011",  "111001110100101111",  "111001110101010011",  "111001110101111000",  "111001110110011100",  "111001110111000001",  "111001110111100110",  "111001111000001011",  "111001111000110001",  "111001111001010110",  "111001111001111100",  "111001111010100010",  "111001111011001000",  "111001111011101110",  "111001111100010101",  "111001111100111011",  "111001111101100010",  "111001111110001001",  "111001111110110001",  "111001111111011000",  "111010000000000000",  "111010000000100111",  "111010000001001111",  "111010000001110111",  "111010000010100000",  "111010000011001000",  "111010000011110001",  "111010000100011010",  "111010000101000011",  "111010000101101100",  "111010000110010110",  "111010000110111111",  "111010000111101001",  "111010001000010011",  "111010001000111101",  "111010001001100111",  "111010001010010010",  "111010001010111100",  "111010001011100111",  "111010001100010010",  "111010001100111101",  "111010001101101000",  "111010001110010100",  "111010001111000000",  "111010001111101011",  "111010010000010111",  "111010010001000100",  "111010010001110000",  "111010010010011100",  "111010010011001001",  "111010010011110110",  "111010010100100011",  "111010010101010000",  "111010010101111101",  "111010010110101011",  "111010010111011000",  "111010011000000110",  "111010011000110100",  "111010011001100010",  "111010011010010001",  "111010011010111111",  "111010011011101110",  "111010011100011100",  "111010011101001011",  "111010011101111010",  "111010011110101010",  "111010011111011001",  "111010100000001001",  "111010100000111000",  "111010100001101000",  "111010100010011000",  "111010100011001000",  "111010100011111001",  "111010100100101001",  "111010100101011010",  "111010100110001010",  "111010100110111011",  "111010100111101100",  "111010101000011110",  "111010101001001111",  "111010101010000000",  "111010101010110010",  "111010101011100100",  "111010101100010110",  "111010101101001000",  "111010101101111010",  "111010101110101101",  "111010101111011111",  "111010110000010010",  "111010110001000101",  "111010110001111000",  "111010110010101011",  "111010110011011110",  "111010110100010001",  "111010110101000101",  "111010110101111000",  "111010110110101100",  "111010110111100000",  "111010111000010100",  "111010111001001000",  "111010111001111101",  "111010111010110001",  "111010111011100110",  "111010111100011010",  "111010111101001111",  "111010111110000100",  "111010111110111001",  "111010111111101111",  "111011000000100100",  "111011000001011010",  "111011000010001111",  "111011000011000101",  "111011000011111011",  "111011000100110001",  "111011000101100111",  "111011000110011101",  "111011000111010100",  "111011001000001010",  "111011001001000001",  "111011001001111000",  "111011001010101111",  "111011001011100110",  "111011001100011101",  "111011001101010100",  "111011001110001100",  "111011001111000011",  "111011001111111011",  "111011010000110010",  "111011010001101010",  "111011010010100010",  "111011010011011010",  "111011010100010011",  "111011010101001011",  "111011010110000011",  "111011010110111100",  "111011010111110101",  "111011011000101101",  "111011011001100110",  "111011011010011111",  "111011011011011000",  "111011011100010010",  "111011011101001011",  "111011011110000100",  "111011011110111110",  "111011011111111000",  "111011100000110001",  "111011100001101011",  "111011100010100101",  "111011100011011111",  "111011100100011001",  "111011100101010100",  "111011100110001110",  "111011100111001001",  "111011101000000011",  "111011101000111110",  "111011101001111001",  "111011101010110100",  "111011101011101111",  "111011101100101010",  "111011101101100101",  "111011101110100000",  "111011101111011100",  "111011110000010111",  "111011110001010011",  "111011110010001110",  "111011110011001010",  "111011110100000110",  "111011110101000010",  "111011110101111110",  "111011110110111010",  "111011110111110110",  "111011111000110011",  "111011111001101111",  "111011111010101100",  "111011111011101000",  "111011111100100101",  "111011111101100010",  "111011111110011111",  "111011111111011100",  "111100000000011001",  "111100000001010110",  "111100000010010011",  "111100000011010000",  "111100000100001110",  "111100000101001011",  "111100000110001000",  "111100000111000110",  "111100001000000100",  "111100001001000010",  "111100001001111111",  "111100001010111101",  "111100001011111011",  "111100001100111001",  "111100001101111000",  "111100001110110110",  "111100001111110100",  "111100010000110010",  "111100010001110001",  "111100010010101111",  "111100010011101110",  "111100010100101101",  "111100010101101100",  "111100010110101010",  "111100010111101001",  "111100011000101000",  "111100011001100111",  "111100011010100110",  "111100011011100101",  "111100011100100101",  "111100011101100100",  "111100011110100011",  "111100011111100011",  "111100100000100010",  "111100100001100010",  "111100100010100001",  "111100100011100001",  "111100100100100001",  "111100100101100001",  "111100100110100001",  "111100100111100000",  "111100101000100000",  "111100101001100000",  "111100101010100001",  "111100101011100001",  "111100101100100001",  "111100101101100001",  "111100101110100010",  "111100101111100010",  "111100110000100010",  "111100110001100011",  "111100110010100011",  "111100110011100100",  "111100110100100101",  "111100110101100101",  "111100110110100110",  "111100110111100111",  "111100111000101000",  "111100111001101001",  "111100111010101010",  "111100111011101011",  "111100111100101100",  "111100111101101101",  "111100111110101110",  "111100111111101111",  "111101000000110000",  "111101000001110001",  "111101000010110011",  "111101000011110100",  "111101000100110101",  "111101000101110111",  "111101000110111000",  "111101000111111010",  "111101001000111011",  "111101001001111101",  "111101001010111111",  "111101001100000000",  "111101001101000010",  "111101001110000100",  "111101001111000110",  "111101010000000111",  "111101010001001001",  "111101010010001011",  "111101010011001101",  "111101010100001111",  "111101010101010001",  "111101010110010011",  "111101010111010101",  "111101011000010111",  "111101011001011001",  "111101011010011011",  "111101011011011101",  "111101011100100000",  "111101011101100010",  "111101011110100100",  "111101011111100110",  "111101100000101001",  "111101100001101011",  "111101100010101101",  "111101100011110000",  "111101100100110010",  "111101100101110100",  "111101100110110111",  "111101100111111001",  "111101101000111100",  "111101101001111110",  "111101101011000001",  "111101101100000011",  "111101101101000110",  "111101101110001000",  "111101101111001011",  "111101110000001101",  "111101110001010000",  "111101110010010011",  "111101110011010101",  "111101110100011000",  "111101110101011010",  "111101110110011101",  "111101110111100000",  "111101111000100010",  "111101111001100101",  "111101111010101000",  "111101111011101011",  "111101111100101101",  "111101111101110000",  "111101111110110011",  "111101111111110110",  "111110000000111000",  "111110000001111011",  "111110000010111110",  "111110000100000001",  "111110000101000011",  "111110000110000110",  "111110000111001001",  "111110001000001100",  "111110001001001110",  "111110001010010001",  "111110001011010100",  "111110001100010111",  "111110001101011010",  "111110001110011100",  "111110001111011111",  "111110010000100010",  "111110010001100101",  "111110010010100111",  "111110010011101010",  "111110010100101101",  "111110010101110000",  "111110010110110010",  "111110010111110101",  "111110011000111000",  "111110011001111011",  "111110011010111101",  "111110011100000000",  "111110011101000011",  "111110011110000101",  "111110011111001000",  "111110100000001011",  "111110100001001101",  "111110100010010000",  "111110100011010011",  "111110100100010101",  "111110100101011000",  "111110100110011010",  "111110100111011101",  "111110101000100000",  "111110101001100010",  "111110101010100101",  "111110101011100111",  "111110101100101010",  "111110101101101100",  "111110101110101110",  "111110101111110001",  "111110110000110011",  "111110110001110110",  "111110110010111000",  "111110110011111010",  "111110110100111101",  "111110110101111111",  "111110110111000001",  "111110111000000011",  "111110111001000110",  "111110111010001000",  "111110111011001010",  "111110111100001100",  "111110111101001110",  "111110111110010000",  "111110111111010010",  "111111000000010100",  "111111000001010110",  "111111000010011000",  "111111000011011010",  "111111000100011100",  "111111000101011110",  "111111000110100000",  "111111000111100010",  "111111001000100011",  "111111001001100101",  "111111001010100111",  "111111001011101000",  "111111001100101010",  "111111001101101100",  "111111001110101101",  "111111001111101111",  "111111010000110000",  "111111010001110001",  "111111010010110011",  "111111010011110100",  "111111010100110110",  "111111010101110111",  "111111010110111000",  "111111010111111001",  "111111011000111010",  "111111011001111011",  "111111011010111100",  "111111011011111110",  "111111011100111110",  "111111011101111111",  "111111011111000000",  "111111100000000001",  "111111100001000010",  "111111100010000011",  "111111100011000011",  "111111100100000100",  "111111100101000101",  "111111100110000101",  "111111100111000110",  "111111101000000110",  "111111101001000110",  "111111101010000111",  "111111101011000111",  "111111101100000111",  "111111101101000111",  "111111101110001000",  "111111101111001000",  "111111110000001000",  "111111110001001000",  "111111110010000111",  "111111110011000111",  "111111110100000111",  "111111110101000111",  "111111110110000111",  "111111110111000110",  "111111111000000110",  "111111111001000101",  "111111111010000101",  "111111111011000100",  "111111111100000011",  "111111111101000011",  "111111111110000010",  "111111111111000001"),("000000000000000000",  "000000000000111111",  "000000000001111110",  "000000000010111101",  "000000000011111100",  "000000000100111010",  "000000000101111001",  "000000000110111000",  "000000000111110110",  "000000001000110101",  "000000001001110011",  "000000001010110001",  "000000001011110000",  "000000001100101110",  "000000001101101100",  "000000001110101010",  "000000001111101000",  "000000010000100110",  "000000010001100100",  "000000010010100010",  "000000010011011111",  "000000010100011101",  "000000010101011011",  "000000010110011000",  "000000010111010101",  "000000011000010011",  "000000011001010000",  "000000011010001101",  "000000011011001010",  "000000011100000111",  "000000011101000100",  "000000011110000001",  "000000011110111110",  "000000011111111011",  "000000100000110111",  "000000100001110100",  "000000100010110000",  "000000100011101101",  "000000100100101001",  "000000100101100101",  "000000100110100010",  "000000100111011110",  "000000101000011010",  "000000101001010101",  "000000101010010001",  "000000101011001101",  "000000101100001001",  "000000101101000100",  "000000101110000000",  "000000101110111011",  "000000101111110110",  "000000110000110010",  "000000110001101101",  "000000110010101000",  "000000110011100011",  "000000110100011110",  "000000110101011000",  "000000110110010011",  "000000110111001110",  "000000111000001000",  "000000111001000011",  "000000111001111101",  "000000111010110111",  "000000111011110001",  "000000111100101011",  "000000111101100101",  "000000111110011111",  "000000111111011001",  "000001000000010011",  "000001000001001100",  "000001000010000110",  "000001000010111111",  "000001000011111000",  "000001000100110001",  "000001000101101011",  "000001000110100100",  "000001000111011100",  "000001001000010101",  "000001001001001110",  "000001001010000111",  "000001001010111111",  "000001001011110111",  "000001001100110000",  "000001001101101000",  "000001001110100000",  "000001001111011000",  "000001010000010000",  "000001010001001000",  "000001010001111111",  "000001010010110111",  "000001010011101110",  "000001010100100110",  "000001010101011101",  "000001010110010100",  "000001010111001011",  "000001011000000010",  "000001011000111001",  "000001011001110000",  "000001011010100111",  "000001011011011101",  "000001011100010011",  "000001011101001010",  "000001011110000000",  "000001011110110110",  "000001011111101100",  "000001100000100010",  "000001100001011000",  "000001100010001101",  "000001100011000011",  "000001100011111000",  "000001100100101110",  "000001100101100011",  "000001100110011000",  "000001100111001101",  "000001101000000010",  "000001101000110111",  "000001101001101011",  "000001101010100000",  "000001101011010100",  "000001101100001001",  "000001101100111101",  "000001101101110001",  "000001101110100101",  "000001101111011001",  "000001110000001100",  "000001110001000000",  "000001110001110011",  "000001110010100111",  "000001110011011010",  "000001110100001101",  "000001110101000000",  "000001110101110011",  "000001110110100110",  "000001110111011001",  "000001111000001011",  "000001111000111101",  "000001111001110000",  "000001111010100010",  "000001111011010100",  "000001111100000110",  "000001111100111000",  "000001111101101001",  "000001111110011011",  "000001111111001100",  "000001111111111110",  "000010000000101111",  "000010000001100000",  "000010000010010001",  "000010000011000010",  "000010000011110011",  "000010000100100011",  "000010000101010100",  "000010000110000100",  "000010000110110100",  "000010000111100100",  "000010001000010100",  "000010001001000100",  "000010001001110100",  "000010001010100011",  "000010001011010011",  "000010001100000010",  "000010001100110001",  "000010001101100000",  "000010001110001111",  "000010001110111110",  "000010001111101100",  "000010010000011011",  "000010010001001001",  "000010010001111000",  "000010010010100110",  "000010010011010100",  "000010010100000010",  "000010010100101111",  "000010010101011101",  "000010010110001010",  "000010010110111000",  "000010010111100101",  "000010011000010010",  "000010011000111111",  "000010011001101100",  "000010011010011000",  "000010011011000101",  "000010011011110001",  "000010011100011110",  "000010011101001010",  "000010011101110110",  "000010011110100010",  "000010011111001101",  "000010011111111001",  "000010100000100100",  "000010100001010000",  "000010100001111011",  "000010100010100110",  "000010100011010001",  "000010100011111100",  "000010100100100110",  "000010100101010001",  "000010100101111011",  "000010100110100101",  "000010100111001111",  "000010100111111001",  "000010101000100011",  "000010101001001101",  "000010101001110110",  "000010101010011111",  "000010101011001001",  "000010101011110010",  "000010101100011011",  "000010101101000011",  "000010101101101100",  "000010101110010101",  "000010101110111101",  "000010101111100101",  "000010110000001101",  "000010110000110101",  "000010110001011101",  "000010110010000101",  "000010110010101100",  "000010110011010100",  "000010110011111011",  "000010110100100010",  "000010110101001001",  "000010110101110000",  "000010110110010110",  "000010110110111101",  "000010110111100011",  "000010111000001001",  "000010111000101111",  "000010111001010101",  "000010111001111011",  "000010111010100001",  "000010111011000110",  "000010111011101011",  "000010111100010001",  "000010111100110110",  "000010111101011011",  "000010111101111111",  "000010111110100100",  "000010111111001000",  "000010111111101101",  "000011000000010001",  "000011000000110101",  "000011000001011001",  "000011000001111100",  "000011000010100000",  "000011000011000011",  "000011000011100110",  "000011000100001010",  "000011000100101101",  "000011000101001111",  "000011000101110010",  "000011000110010100",  "000011000110110111",  "000011000111011001",  "000011000111111011",  "000011001000011101",  "000011001000111111",  "000011001001100000",  "000011001010000010",  "000011001010100011",  "000011001011000100",  "000011001011100101",  "000011001100000110",  "000011001100100111",  "000011001101000111",  "000011001101101000",  "000011001110001000",  "000011001110101000",  "000011001111001000",  "000011001111100111",  "000011010000000111",  "000011010000100111",  "000011010001000110",  "000011010001100101",  "000011010010000100",  "000011010010100011",  "000011010011000001",  "000011010011100000",  "000011010011111110",  "000011010100011101",  "000011010100111011",  "000011010101011001",  "000011010101110110",  "000011010110010100",  "000011010110110001",  "000011010111001111",  "000011010111101100",  "000011011000001001",  "000011011000100101",  "000011011001000010",  "000011011001011111",  "000011011001111011",  "000011011010010111",  "000011011010110011",  "000011011011001111",  "000011011011101011",  "000011011100000110",  "000011011100100010",  "000011011100111101",  "000011011101011000",  "000011011101110011",  "000011011110001110",  "000011011110101000",  "000011011111000011",  "000011011111011101",  "000011011111110111",  "000011100000010001",  "000011100000101011",  "000011100001000101",  "000011100001011110",  "000011100001111000",  "000011100010010001",  "000011100010101010",  "000011100011000011",  "000011100011011011",  "000011100011110100",  "000011100100001100",  "000011100100100100",  "000011100100111101",  "000011100101010100",  "000011100101101100",  "000011100110000100",  "000011100110011011",  "000011100110110011",  "000011100111001010",  "000011100111100001",  "000011100111110111",  "000011101000001110",  "000011101000100101",  "000011101000111011",  "000011101001010001",  "000011101001100111",  "000011101001111101",  "000011101010010010",  "000011101010101000",  "000011101010111101",  "000011101011010011",  "000011101011101000",  "000011101011111100",  "000011101100010001",  "000011101100100110",  "000011101100111010",  "000011101101001110",  "000011101101100010",  "000011101101110110",  "000011101110001010",  "000011101110011110",  "000011101110110001",  "000011101111000100",  "000011101111010111",  "000011101111101010",  "000011101111111101",  "000011110000010000",  "000011110000100010",  "000011110000110101",  "000011110001000111",  "000011110001011001",  "000011110001101010",  "000011110001111100",  "000011110010001110",  "000011110010011111",  "000011110010110000",  "000011110011000001",  "000011110011010010",  "000011110011100011",  "000011110011110011",  "000011110100000100",  "000011110100010100",  "000011110100100100",  "000011110100110100",  "000011110101000011",  "000011110101010011",  "000011110101100010",  "000011110101110010",  "000011110110000001",  "000011110110010000",  "000011110110011110",  "000011110110101101",  "000011110110111011",  "000011110111001010",  "000011110111011000",  "000011110111100110",  "000011110111110011",  "000011111000000001",  "000011111000001110",  "000011111000011100",  "000011111000101001",  "000011111000110110",  "000011111001000011",  "000011111001001111",  "000011111001011100",  "000011111001101000",  "000011111001110100",  "000011111010000000",  "000011111010001100",  "000011111010011000",  "000011111010100011",  "000011111010101111",  "000011111010111010",  "000011111011000101",  "000011111011010000",  "000011111011011011",  "000011111011100101",  "000011111011110000",  "000011111011111010",  "000011111100000100",  "000011111100001110",  "000011111100011000",  "000011111100100001",  "000011111100101011",  "000011111100110100",  "000011111100111101",  "000011111101000110",  "000011111101001111",  "000011111101010111",  "000011111101100000",  "000011111101101000",  "000011111101110000",  "000011111101111000",  "000011111110000000",  "000011111110001000",  "000011111110001111",  "000011111110010111",  "000011111110011110",  "000011111110100101",  "000011111110101100",  "000011111110110010",  "000011111110111001",  "000011111110111111",  "000011111111000110",  "000011111111001100",  "000011111111010010",  "000011111111010111",  "000011111111011101",  "000011111111100010",  "000011111111101000",  "000011111111101101",  "000011111111110010",  "000011111111110110",  "000011111111111011",  "000100000000000000",  "000100000000000100",  "000100000000001000",  "000100000000001100",  "000100000000010000",  "000100000000010100",  "000100000000010111",  "000100000000011011",  "000100000000011110",  "000100000000100001",  "000100000000100100",  "000100000000100111",  "000100000000101001",  "000100000000101100",  "000100000000101110",  "000100000000110000",  "000100000000110010",  "000100000000110100",  "000100000000110101",  "000100000000110111",  "000100000000111000",  "000100000000111001",  "000100000000111010",  "000100000000111011",  "000100000000111100",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111101",  "000100000000111100",  "000100000000111011",  "000100000000111011",  "000100000000111010",  "000100000000111001",  "000100000000110111",  "000100000000110110",  "000100000000110100",  "000100000000110010",  "000100000000110000",  "000100000000101110",  "000100000000101100",  "000100000000101010",  "000100000000100111",  "000100000000100101",  "000100000000100010",  "000100000000011111",  "000100000000011100",  "000100000000011000",  "000100000000010101",  "000100000000010001",  "000100000000001110",  "000100000000001010",  "000100000000000110",  "000100000000000001",  "000011111111111101",  "000011111111111001",  "000011111111110100",  "000011111111101111",  "000011111111101010",  "000011111111100101",  "000011111111100000",  "000011111111011010",  "000011111111010101",  "000011111111001111",  "000011111111001001",  "000011111111000011",  "000011111110111101",  "000011111110110111",  "000011111110110000",  "000011111110101010",  "000011111110100011",  "000011111110011100",  "000011111110010101",  "000011111110001110",  "000011111110000111",  "000011111101111111",  "000011111101111000",  "000011111101110000",  "000011111101101000",  "000011111101100000",  "000011111101011000",  "000011111101001111",  "000011111101000111",  "000011111100111110",  "000011111100110101",  "000011111100101100",  "000011111100100011",  "000011111100011010",  "000011111100010001",  "000011111100000111",  "000011111011111101",  "000011111011110100",  "000011111011101010",  "000011111011100000",  "000011111011010101",  "000011111011001011",  "000011111011000000",  "000011111010110110",  "000011111010101011",  "000011111010100000",  "000011111010010101",  "000011111010001010",  "000011111001111110",  "000011111001110011",  "000011111001100111",  "000011111001011011",  "000011111001001111",  "000011111001000011",  "000011111000110111",  "000011111000101011",  "000011111000011110",  "000011111000010001",  "000011111000000101",  "000011110111111000",  "000011110111101011",  "000011110111011101",  "000011110111010000",  "000011110111000011",  "000011110110110101",  "000011110110100111",  "000011110110011001",  "000011110110001011",  "000011110101111101",  "000011110101101111",  "000011110101100000",  "000011110101010010",  "000011110101000011",  "000011110100110100",  "000011110100100101",  "000011110100010110",  "000011110100000111",  "000011110011110111",  "000011110011101000",  "000011110011011000",  "000011110011001000",  "000011110010111000",  "000011110010101000",  "000011110010011000",  "000011110010001000",  "000011110001110111",  "000011110001100111",  "000011110001010110",  "000011110001000101",  "000011110000110100",  "000011110000100011",  "000011110000010010",  "000011110000000000",  "000011101111101111",  "000011101111011101",  "000011101111001011",  "000011101110111001",  "000011101110100111",  "000011101110010101",  "000011101110000011",  "000011101101110000",  "000011101101011110",  "000011101101001011",  "000011101100111000",  "000011101100100101",  "000011101100010010",  "000011101011111111",  "000011101011101100",  "000011101011011000",  "000011101011000101",  "000011101010110001",  "000011101010011101",  "000011101010001001",  "000011101001110101",  "000011101001100001",  "000011101001001101",  "000011101000111000",  "000011101000100011",  "000011101000001111",  "000011100111111010",  "000011100111100101",  "000011100111010000",  "000011100110111011",  "000011100110100101",  "000011100110010000",  "000011100101111010",  "000011100101100101",  "000011100101001111",  "000011100100111001",  "000011100100100011",  "000011100100001101",  "000011100011110110",  "000011100011100000",  "000011100011001001",  "000011100010110011",  "000011100010011100",  "000011100010000101",  "000011100001101110",  "000011100001010111",  "000011100001000000",  "000011100000101000",  "000011100000010001",  "000011011111111001",  "000011011111100001",  "000011011111001010",  "000011011110110010",  "000011011110011010",  "000011011110000001",  "000011011101101001",  "000011011101010001",  "000011011100111000",  "000011011100011111",  "000011011100000111",  "000011011011101110",  "000011011011010101",  "000011011010111100",  "000011011010100011",  "000011011010001001",  "000011011001110000",  "000011011001010110",  "000011011000111101",  "000011011000100011",  "000011011000001001",  "000011010111101111",  "000011010111010101",  "000011010110111011",  "000011010110100000",  "000011010110000110",  "000011010101101011",  "000011010101010001",  "000011010100110110",  "000011010100011011",  "000011010100000000",  "000011010011100101",  "000011010011001010",  "000011010010101111",  "000011010010010011",  "000011010001111000",  "000011010001011100",  "000011010001000000",  "000011010000100101",  "000011010000001001",  "000011001111101101",  "000011001111010000",  "000011001110110100",  "000011001110011000",  "000011001101111011",  "000011001101011111",  "000011001101000010",  "000011001100100110",  "000011001100001001",  "000011001011101100",  "000011001011001111",  "000011001010110010",  "000011001010010100",  "000011001001110111",  "000011001001011010",  "000011001000111100",  "000011001000011110",  "000011001000000001",  "000011000111100011",  "000011000111000101",  "000011000110100111",  "000011000110001001",  "000011000101101010",  "000011000101001100",  "000011000100101110",  "000011000100001111",  "000011000011110001",  "000011000011010010",  "000011000010110011",  "000011000010010100",  "000011000001110101",  "000011000001010110",  "000011000000110111",  "000011000000011000",  "000010111111111000",  "000010111111011001",  "000010111110111001",  "000010111110011010",  "000010111101111010",  "000010111101011010",  "000010111100111010",  "000010111100011010",  "000010111011111010",  "000010111011011010",  "000010111010111010",  "000010111010011001",  "000010111001111001",  "000010111001011001",  "000010111000111000",  "000010111000010111",  "000010110111110110",  "000010110111010110",  "000010110110110101",  "000010110110010100",  "000010110101110010",  "000010110101010001",  "000010110100110000",  "000010110100001111",  "000010110011101101",  "000010110011001100",  "000010110010101010",  "000010110010001000",  "000010110001100110",  "000010110001000101",  "000010110000100011",  "000010110000000001",  "000010101111011110",  "000010101110111100",  "000010101110011010",  "000010101101111000",  "000010101101010101",  "000010101100110011",  "000010101100010000",  "000010101011101101",  "000010101011001011",  "000010101010101000",  "000010101010000101",  "000010101001100010",  "000010101000111111",  "000010101000011100",  "000010100111111001",  "000010100111010101",  "000010100110110010",  "000010100110001111",  "000010100101101011",  "000010100101001000",  "000010100100100100",  "000010100100000000",  "000010100011011100",  "000010100010111001",  "000010100010010101",  "000010100001110001",  "000010100001001101",  "000010100000101000",  "000010100000000100",  "000010011111100000",  "000010011110111100",  "000010011110010111",  "000010011101110011",  "000010011101001110",  "000010011100101001",  "000010011100000101",  "000010011011100000",  "000010011010111011",  "000010011010010110",  "000010011001110001",  "000010011001001100",  "000010011000100111",  "000010011000000010",  "000010010111011101",  "000010010110111000",  "000010010110010010",  "000010010101101101",  "000010010101000111",  "000010010100100010",  "000010010011111100",  "000010010011010111",  "000010010010110001",  "000010010010001011",  "000010010001100101",  "000010010000111111",  "000010010000011001",  "000010001111110011",  "000010001111001101",  "000010001110100111",  "000010001110000001",  "000010001101011011",  "000010001100110100",  "000010001100001110",  "000010001011101000",  "000010001011000001",  "000010001010011011",  "000010001001110100",  "000010001001001101",  "000010001000100111",  "000010001000000000",  "000010000111011001",  "000010000110110010",  "000010000110001011",  "000010000101100101",  "000010000100111110",  "000010000100010110",  "000010000011101111",  "000010000011001000",  "000010000010100001",  "000010000001111010",  "000010000001010010",  "000010000000101011",  "000010000000000100",  "000001111111011100",  "000001111110110101",  "000001111110001101",  "000001111101100110",  "000001111100111110",  "000001111100010110",  "000001111011101110",  "000001111011000111",  "000001111010011111",  "000001111001110111",  "000001111001001111",  "000001111000100111",  "000001110111111111",  "000001110111010111",  "000001110110101111",  "000001110110000111",  "000001110101011111",  "000001110100110110",  "000001110100001110",  "000001110011100110",  "000001110010111110",  "000001110010010101",  "000001110001101101",  "000001110001000100",  "000001110000011100",  "000001101111110011",  "000001101111001011",  "000001101110100010",  "000001101101111001",  "000001101101010001",  "000001101100101000",  "000001101011111111",  "000001101011010111",  "000001101010101110",  "000001101010000101",  "000001101001011100",  "000001101000110011",  "000001101000001010",  "000001100111100001",  "000001100110111000",  "000001100110001111",  "000001100101100110",  "000001100100111101",  "000001100100010100",  "000001100011101010",  "000001100011000001",  "000001100010011000",  "000001100001101111",  "000001100001000101",  "000001100000011100",  "000001011111110011",  "000001011111001001",  "000001011110100000",  "000001011101110111",  "000001011101001101",  "000001011100100100",  "000001011011111010",  "000001011011010001",  "000001011010100111",  "000001011001111101",  "000001011001010100",  "000001011000101010",  "000001011000000000",  "000001010111010111",  "000001010110101101",  "000001010110000011",  "000001010101011010",  "000001010100110000",  "000001010100000110",  "000001010011011100",  "000001010010110010",  "000001010010001000",  "000001010001011111",  "000001010000110101",  "000001010000001011",  "000001001111100001",  "000001001110110111",  "000001001110001101",  "000001001101100011",  "000001001100111001",  "000001001100001111",  "000001001011100101",  "000001001010111011",  "000001001010010001",  "000001001001100111",  "000001001000111101",  "000001001000010011",  "000001000111101000",  "000001000110111110",  "000001000110010100",  "000001000101101010",  "000001000101000000",  "000001000100010110",  "000001000011101011",  "000001000011000001",  "000001000010010111",  "000001000001101101",  "000001000001000011",  "000001000000011000",  "000000111111101110",  "000000111111000100",  "000000111110011010",  "000000111101101111",  "000000111101000101",  "000000111100011011",  "000000111011110000",  "000000111011000110",  "000000111010011100",  "000000111001110010",  "000000111001000111",  "000000111000011101",  "000000110111110011",  "000000110111001000",  "000000110110011110",  "000000110101110100",  "000000110101001001",  "000000110100011111",  "000000110011110101",  "000000110011001010",  "000000110010100000",  "000000110001110110",  "000000110001001011",  "000000110000100001",  "000000101111110111",  "000000101111001100",  "000000101110100010",  "000000101101111000",  "000000101101001101",  "000000101100100011",  "000000101011111001",  "000000101011001110",  "000000101010100100",  "000000101001111010",  "000000101001001111",  "000000101000100101",  "000000100111111011",  "000000100111010000",  "000000100110100110",  "000000100101111100",  "000000100101010010",  "000000100100100111",  "000000100011111101",  "000000100011010011",  "000000100010101001",  "000000100001111110",  "000000100001010100",  "000000100000101010",  "000000100000000000",  "000000011111010110",  "000000011110101011",  "000000011110000001",  "000000011101010111",  "000000011100101101",  "000000011100000011",  "000000011011011001",  "000000011010101111",  "000000011010000100",  "000000011001011010",  "000000011000110000",  "000000011000000110",  "000000010111011100",  "000000010110110010",  "000000010110001000",  "000000010101011110",  "000000010100110100",  "000000010100001010",  "000000010011100000",  "000000010010110110",  "000000010010001100",  "000000010001100011",  "000000010000111001",  "000000010000001111",  "000000001111100101",  "000000001110111011",  "000000001110010001",  "000000001101101000",  "000000001100111110",  "000000001100010100",  "000000001011101011",  "000000001011000001",  "000000001010010111",  "000000001001101110",  "000000001001000100",  "000000001000011010",  "000000000111110001",  "000000000111000111",  "000000000110011110",  "000000000101110100",  "000000000101001011",  "000000000100100001",  "000000000011111000",  "000000000011001111",  "000000000010100101",  "000000000001111100",  "000000000001010011",  "000000000000101001"),("000000000000000000",  "111111111111010111",  "111111111110101110",  "111111111110000100",  "111111111101011011",  "111111111100110010",  "111111111100001001",  "111111111011100000",  "111111111010110111",  "111111111010001110",  "111111111001100101",  "111111111000111100",  "111111111000010011",  "111111110111101011",  "111111110111000010",  "111111110110011001",  "111111110101110000",  "111111110101000111",  "111111110100011111",  "111111110011110110",  "111111110011001110",  "111111110010100101",  "111111110001111100",  "111111110001010100",  "111111110000101011",  "111111110000000011",  "111111101111011011",  "111111101110110010",  "111111101110001010",  "111111101101100010",  "111111101100111001",  "111111101100010001",  "111111101011101001",  "111111101011000001",  "111111101010011001",  "111111101001110001",  "111111101001001001",  "111111101000100001",  "111111100111111001",  "111111100111010001",  "111111100110101001",  "111111100110000010",  "111111100101011010",  "111111100100110010",  "111111100100001011",  "111111100011100011",  "111111100010111011",  "111111100010010100",  "111111100001101100",  "111111100001000101",  "111111100000011110",  "111111011111110110",  "111111011111001111",  "111111011110101000",  "111111011110000000",  "111111011101011001",  "111111011100110010",  "111111011100001011",  "111111011011100100",  "111111011010111101",  "111111011010010110",  "111111011001101111",  "111111011001001001",  "111111011000100010",  "111111010111111011",  "111111010111010100",  "111111010110101110",  "111111010110000111",  "111111010101100001",  "111111010100111010",  "111111010100010100",  "111111010011101110",  "111111010011000111",  "111111010010100001",  "111111010001111011",  "111111010001010101",  "111111010000101111",  "111111010000001001",  "111111001111100011",  "111111001110111101",  "111111001110010111",  "111111001101110001",  "111111001101001011",  "111111001100100110",  "111111001100000000",  "111111001011011010",  "111111001010110101",  "111111001010001111",  "111111001001101010",  "111111001001000101",  "111111001000011111",  "111111000111111010",  "111111000111010101",  "111111000110110000",  "111111000110001011",  "111111000101100110",  "111111000101000001",  "111111000100011100",  "111111000011110111",  "111111000011010011",  "111111000010101110",  "111111000010001001",  "111111000001100101",  "111111000001000000",  "111111000000011100",  "111110111111110111",  "111110111111010011",  "111110111110101111",  "111110111110001011",  "111110111101100110",  "111110111101000010",  "111110111100011110",  "111110111011111010",  "111110111011010111",  "111110111010110011",  "111110111010001111",  "111110111001101011",  "111110111001001000",  "111110111000100100",  "111110111000000001",  "111110110111011101",  "111110110110111010",  "111110110110010111",  "111110110101110100",  "111110110101010001",  "111110110100101110",  "111110110100001011",  "111110110011101000",  "111110110011000101",  "111110110010100010",  "111110110001111111",  "111110110001011101",  "111110110000111010",  "111110110000011000",  "111110101111110101",  "111110101111010011",  "111110101110110001",  "111110101110001110",  "111110101101101100",  "111110101101001010",  "111110101100101000",  "111110101100000110",  "111110101011100100",  "111110101011000011",  "111110101010100001",  "111110101001111111",  "111110101001011110",  "111110101000111100",  "111110101000011011",  "111110100111111010",  "111110100111011000",  "111110100110110111",  "111110100110010110",  "111110100101110101",  "111110100101010100",  "111110100100110011",  "111110100100010010",  "111110100011110010",  "111110100011010001",  "111110100010110000",  "111110100010010000",  "111110100001110000",  "111110100001001111",  "111110100000101111",  "111110100000001111",  "111110011111101111",  "111110011111001111",  "111110011110101111",  "111110011110001111",  "111110011101101111",  "111110011101010000",  "111110011100110000",  "111110011100010000",  "111110011011110001",  "111110011011010010",  "111110011010110010",  "111110011010010011",  "111110011001110100",  "111110011001010101",  "111110011000110110",  "111110011000010111",  "111110010111111000",  "111110010111011010",  "111110010110111011",  "111110010110011100",  "111110010101111110",  "111110010101100000",  "111110010101000001",  "111110010100100011",  "111110010100000101",  "111110010011100111",  "111110010011001001",  "111110010010101011",  "111110010010001101",  "111110010001110000",  "111110010001010010",  "111110010000110101",  "111110010000010111",  "111110001111111010",  "111110001111011101",  "111110001110111111",  "111110001110100010",  "111110001110000101",  "111110001101101000",  "111110001101001100",  "111110001100101111",  "111110001100010010",  "111110001011110110",  "111110001011011001",  "111110001010111101",  "111110001010100001",  "111110001010000100",  "111110001001101000",  "111110001001001100",  "111110001000110000",  "111110001000010101",  "111110000111111001",  "111110000111011101",  "111110000111000010",  "111110000110100110",  "111110000110001011",  "111110000101101111",  "111110000101010100",  "111110000100111001",  "111110000100011110",  "111110000100000011",  "111110000011101000",  "111110000011001110",  "111110000010110011",  "111110000010011000",  "111110000001111110",  "111110000001100100",  "111110000001001001",  "111110000000101111",  "111110000000010101",  "111101111111111011",  "111101111111100001",  "111101111111000111",  "111101111110101110",  "111101111110010100",  "111101111101111011",  "111101111101100001",  "111101111101001000",  "111101111100101111",  "111101111100010110",  "111101111011111100",  "111101111011100100",  "111101111011001011",  "111101111010110010",  "111101111010011001",  "111101111010000001",  "111101111001101000",  "111101111001010000",  "111101111000111000",  "111101111000011111",  "111101111000000111",  "111101110111101111",  "111101110111011000",  "111101110111000000",  "111101110110101000",  "111101110110010001",  "111101110101111001",  "111101110101100010",  "111101110101001010",  "111101110100110011",  "111101110100011100",  "111101110100000101",  "111101110011101110",  "111101110011010111",  "111101110011000001",  "111101110010101010",  "111101110010010100",  "111101110001111101",  "111101110001100111",  "111101110001010001",  "111101110000111011",  "111101110000100101",  "111101110000001111",  "111101101111111001",  "111101101111100011",  "111101101111001110",  "111101101110111000",  "111101101110100011",  "111101101110001110",  "111101101101111000",  "111101101101100011",  "111101101101001110",  "111101101100111010",  "111101101100100101",  "111101101100010000",  "111101101011111100",  "111101101011100111",  "111101101011010011",  "111101101010111111",  "111101101010101010",  "111101101010010110",  "111101101010000010",  "111101101001101111",  "111101101001011011",  "111101101001000111",  "111101101000110100",  "111101101000100000",  "111101101000001101",  "111101100111111010",  "111101100111100111",  "111101100111010100",  "111101100111000001",  "111101100110101110",  "111101100110011011",  "111101100110001001",  "111101100101110110",  "111101100101100100",  "111101100101010001",  "111101100100111111",  "111101100100101101",  "111101100100011011",  "111101100100001001",  "111101100011111000",  "111101100011100110",  "111101100011010100",  "111101100011000011",  "111101100010110010",  "111101100010100000",  "111101100010001111",  "111101100001111110",  "111101100001101101",  "111101100001011101",  "111101100001001100",  "111101100000111011",  "111101100000101011",  "111101100000011010",  "111101100000001010",  "111101011111111010",  "111101011111101010",  "111101011111011010",  "111101011111001010",  "111101011110111010",  "111101011110101011",  "111101011110011011",  "111101011110001100",  "111101011101111101",  "111101011101101101",  "111101011101011110",  "111101011101001111",  "111101011101000000",  "111101011100110010",  "111101011100100011",  "111101011100010100",  "111101011100000110",  "111101011011111000",  "111101011011101001",  "111101011011011011",  "111101011011001101",  "111101011010111111",  "111101011010110010",  "111101011010100100",  "111101011010010110",  "111101011010001001",  "111101011001111100",  "111101011001101110",  "111101011001100001",  "111101011001010100",  "111101011001000111",  "111101011000111010",  "111101011000101110",  "111101011000100001",  "111101011000010101",  "111101011000001000",  "111101010111111100",  "111101010111110000",  "111101010111100100",  "111101010111011000",  "111101010111001100",  "111101010111000000",  "111101010110110101",  "111101010110101001",  "111101010110011110",  "111101010110010011",  "111101010110000111",  "111101010101111100",  "111101010101110001",  "111101010101100111",  "111101010101011100",  "111101010101010001",  "111101010101000111",  "111101010100111100",  "111101010100110010",  "111101010100101000",  "111101010100011110",  "111101010100010100",  "111101010100001010",  "111101010100000000",  "111101010011110110",  "111101010011101101",  "111101010011100100",  "111101010011011010",  "111101010011010001",  "111101010011001000",  "111101010010111111",  "111101010010110110",  "111101010010101101",  "111101010010100101",  "111101010010011100",  "111101010010010100",  "111101010010001011",  "111101010010000011",  "111101010001111011",  "111101010001110011",  "111101010001101011",  "111101010001100100",  "111101010001011100",  "111101010001010100",  "111101010001001101",  "111101010001000110",  "111101010000111110",  "111101010000110111",  "111101010000110000",  "111101010000101001",  "111101010000100011",  "111101010000011100",  "111101010000010101",  "111101010000001111",  "111101010000001001",  "111101010000000010",  "111101001111111100",  "111101001111110110",  "111101001111110000",  "111101001111101011",  "111101001111100101",  "111101001111011111",  "111101001111011010",  "111101001111010101",  "111101001111001111",  "111101001111001010",  "111101001111000101",  "111101001111000000",  "111101001110111100",  "111101001110110111",  "111101001110110010",  "111101001110101110",  "111101001110101001",  "111101001110100101",  "111101001110100001",  "111101001110011101",  "111101001110011001",  "111101001110010101",  "111101001110010010",  "111101001110001110",  "111101001110001011",  "111101001110000111",  "111101001110000100",  "111101001110000001",  "111101001101111110",  "111101001101111011",  "111101001101111000",  "111101001101110101",  "111101001101110011",  "111101001101110000",  "111101001101101110",  "111101001101101100",  "111101001101101001",  "111101001101100111",  "111101001101100101",  "111101001101100100",  "111101001101100010",  "111101001101100000",  "111101001101011111",  "111101001101011101",  "111101001101011100",  "111101001101011011",  "111101001101011010",  "111101001101011001",  "111101001101011000",  "111101001101010111",  "111101001101010111",  "111101001101010110",  "111101001101010110",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010101",  "111101001101010110",  "111101001101010110",  "111101001101010111",  "111101001101010111",  "111101001101011000",  "111101001101011001",  "111101001101011010",  "111101001101011011",  "111101001101011100",  "111101001101011101",  "111101001101011111",  "111101001101100000",  "111101001101100010",  "111101001101100100",  "111101001101100101",  "111101001101100111",  "111101001101101001",  "111101001101101100",  "111101001101101110",  "111101001101110000",  "111101001101110011",  "111101001101110101",  "111101001101111000",  "111101001101111011",  "111101001101111110",  "111101001110000001",  "111101001110000100",  "111101001110000111",  "111101001110001010",  "111101001110001110",  "111101001110010001",  "111101001110010101",  "111101001110011001",  "111101001110011100",  "111101001110100000",  "111101001110100100",  "111101001110101001",  "111101001110101101",  "111101001110110001",  "111101001110110110",  "111101001110111010",  "111101001110111111",  "111101001111000100",  "111101001111001001",  "111101001111001110",  "111101001111010011",  "111101001111011000",  "111101001111011101",  "111101001111100011",  "111101001111101000",  "111101001111101110",  "111101001111110011",  "111101001111111001",  "111101001111111111",  "111101010000000101",  "111101010000001011",  "111101010000010001",  "111101010000011000",  "111101010000011110",  "111101010000100101",  "111101010000101011",  "111101010000110010",  "111101010000111001",  "111101010001000000",  "111101010001000111",  "111101010001001110",  "111101010001010101",  "111101010001011101",  "111101010001100100",  "111101010001101100",  "111101010001110011",  "111101010001111011",  "111101010010000011",  "111101010010001011",  "111101010010010011",  "111101010010011011",  "111101010010100011",  "111101010010101100",  "111101010010110100",  "111101010010111101",  "111101010011000101",  "111101010011001110",  "111101010011010111",  "111101010011100000",  "111101010011101001",  "111101010011110010",  "111101010011111011",  "111101010100000100",  "111101010100001110",  "111101010100010111",  "111101010100100001",  "111101010100101011",  "111101010100110101",  "111101010100111111",  "111101010101001001",  "111101010101010011",  "111101010101011101",  "111101010101100111",  "111101010101110010",  "111101010101111100",  "111101010110000111",  "111101010110010001",  "111101010110011100",  "111101010110100111",  "111101010110110010",  "111101010110111101",  "111101010111001000",  "111101010111010100",  "111101010111011111",  "111101010111101010",  "111101010111110110",  "111101011000000010",  "111101011000001101",  "111101011000011001",  "111101011000100101",  "111101011000110001",  "111101011000111101",  "111101011001001001",  "111101011001010110",  "111101011001100010",  "111101011001101111",  "111101011001111011",  "111101011010001000",  "111101011010010101",  "111101011010100010",  "111101011010101111",  "111101011010111100",  "111101011011001001",  "111101011011010110",  "111101011011100011",  "111101011011110001",  "111101011011111110",  "111101011100001100",  "111101011100011001",  "111101011100100111",  "111101011100110101",  "111101011101000011",  "111101011101010001",  "111101011101011111",  "111101011101101110",  "111101011101111100",  "111101011110001010",  "111101011110011001",  "111101011110100111",  "111101011110110110",  "111101011111000101",  "111101011111010100",  "111101011111100011",  "111101011111110010",  "111101100000000001",  "111101100000010000",  "111101100000011111",  "111101100000101111",  "111101100000111110",  "111101100001001110",  "111101100001011101",  "111101100001101101",  "111101100001111101",  "111101100010001101",  "111101100010011101",  "111101100010101101",  "111101100010111101",  "111101100011001101",  "111101100011011101",  "111101100011101110",  "111101100011111110",  "111101100100001111",  "111101100100100000",  "111101100100110000",  "111101100101000001",  "111101100101010010",  "111101100101100011",  "111101100101110100",  "111101100110000101",  "111101100110010111",  "111101100110101000",  "111101100110111001",  "111101100111001011",  "111101100111011100",  "111101100111101110",  "111101101000000000",  "111101101000010010",  "111101101000100011",  "111101101000110101",  "111101101001000111",  "111101101001011010",  "111101101001101100",  "111101101001111110",  "111101101010010001",  "111101101010100011",  "111101101010110110",  "111101101011001000",  "111101101011011011",  "111101101011101110",  "111101101100000000",  "111101101100010011",  "111101101100100110",  "111101101100111001",  "111101101101001101",  "111101101101100000",  "111101101101110011",  "111101101110000111",  "111101101110011010",  "111101101110101110",  "111101101111000001",  "111101101111010101",  "111101101111101001",  "111101101111111101",  "111101110000010001",  "111101110000100101",  "111101110000111001",  "111101110001001101",  "111101110001100001",  "111101110001110101",  "111101110010001010",  "111101110010011110",  "111101110010110011",  "111101110011000111",  "111101110011011100",  "111101110011110001",  "111101110100000110",  "111101110100011010",  "111101110100101111",  "111101110101000100",  "111101110101011010",  "111101110101101111",  "111101110110000100",  "111101110110011001",  "111101110110101111",  "111101110111000100",  "111101110111011010",  "111101110111101111",  "111101111000000101",  "111101111000011011",  "111101111000110000",  "111101111001000110",  "111101111001011100",  "111101111001110010",  "111101111010001000",  "111101111010011111",  "111101111010110101",  "111101111011001011",  "111101111011100001",  "111101111011111000",  "111101111100001110",  "111101111100100101",  "111101111100111011",  "111101111101010010",  "111101111101101001",  "111101111110000000",  "111101111110010111",  "111101111110101110",  "111101111111000101",  "111101111111011100",  "111101111111110011",  "111110000000001010",  "111110000000100001",  "111110000000111001",  "111110000001010000",  "111110000001100111",  "111110000001111111",  "111110000010010110",  "111110000010101110",  "111110000011000110",  "111110000011011110",  "111110000011110101",  "111110000100001101",  "111110000100100101",  "111110000100111101",  "111110000101010101",  "111110000101101101",  "111110000110000110",  "111110000110011110",  "111110000110110110",  "111110000111001111",  "111110000111100111",  "111110001000000000",  "111110001000011000",  "111110001000110001",  "111110001001001001",  "111110001001100010",  "111110001001111011",  "111110001010010100",  "111110001010101101",  "111110001011000101",  "111110001011011110",  "111110001011111000",  "111110001100010001",  "111110001100101010",  "111110001101000011",  "111110001101011100",  "111110001101110110",  "111110001110001111",  "111110001110101000",  "111110001111000010",  "111110001111011100",  "111110001111110101",  "111110010000001111",  "111110010000101001",  "111110010001000010",  "111110010001011100",  "111110010001110110",  "111110010010010000",  "111110010010101010",  "111110010011000100",  "111110010011011110",  "111110010011111000",  "111110010100010010",  "111110010100101100",  "111110010101000111",  "111110010101100001",  "111110010101111011",  "111110010110010110",  "111110010110110000",  "111110010111001011",  "111110010111100101",  "111110011000000000",  "111110011000011011",  "111110011000110101",  "111110011001010000",  "111110011001101011",  "111110011010000110",  "111110011010100001",  "111110011010111100",  "111110011011010111",  "111110011011110010",  "111110011100001101",  "111110011100101000",  "111110011101000011",  "111110011101011110",  "111110011101111001",  "111110011110010101",  "111110011110110000",  "111110011111001011",  "111110011111100111",  "111110100000000010",  "111110100000011110",  "111110100000111001",  "111110100001010101",  "111110100001110001",  "111110100010001100",  "111110100010101000",  "111110100011000100",  "111110100011100000",  "111110100011111011",  "111110100100010111",  "111110100100110011",  "111110100101001111",  "111110100101101011",  "111110100110000111",  "111110100110100011",  "111110100110111111",  "111110100111011011",  "111110100111111000",  "111110101000010100",  "111110101000110000",  "111110101001001100",  "111110101001101001",  "111110101010000101",  "111110101010100010",  "111110101010111110",  "111110101011011010",  "111110101011110111",  "111110101100010011",  "111110101100110000",  "111110101101001101",  "111110101101101001",  "111110101110000110",  "111110101110100011",  "111110101110111111",  "111110101111011100",  "111110101111111001",  "111110110000010110",  "111110110000110011",  "111110110001010000",  "111110110001101101",  "111110110010001010",  "111110110010100111",  "111110110011000100",  "111110110011100001",  "111110110011111110",  "111110110100011011",  "111110110100111000",  "111110110101010101",  "111110110101110010",  "111110110110010000",  "111110110110101101",  "111110110111001010",  "111110110111100111",  "111110111000000101",  "111110111000100010",  "111110111001000000",  "111110111001011101",  "111110111001111010",  "111110111010011000",  "111110111010110101",  "111110111011010011",  "111110111011110000",  "111110111100001110",  "111110111100101100",  "111110111101001001",  "111110111101100111",  "111110111110000101",  "111110111110100010",  "111110111111000000",  "111110111111011110",  "111110111111111100",  "111111000000011001",  "111111000000110111",  "111111000001010101",  "111111000001110011",  "111111000010010001",  "111111000010101111",  "111111000011001100",  "111111000011101010",  "111111000100001000",  "111111000100100110",  "111111000101000100",  "111111000101100010",  "111111000110000000",  "111111000110011110",  "111111000110111100",  "111111000111011010",  "111111000111111001",  "111111001000010111",  "111111001000110101",  "111111001001010011",  "111111001001110001",  "111111001010001111",  "111111001010101101",  "111111001011001100",  "111111001011101010",  "111111001100001000",  "111111001100100110",  "111111001101000101",  "111111001101100011",  "111111001110000001",  "111111001110100000",  "111111001110111110",  "111111001111011100",  "111111001111111010",  "111111010000011001",  "111111010000110111",  "111111010001010110",  "111111010001110100",  "111111010010010010",  "111111010010110001",  "111111010011001111",  "111111010011101110",  "111111010100001100",  "111111010100101011",  "111111010101001001",  "111111010101100111",  "111111010110000110",  "111111010110100100",  "111111010111000011",  "111111010111100001",  "111111011000000000",  "111111011000011110",  "111111011000111101",  "111111011001011011",  "111111011001111010",  "111111011010011001",  "111111011010110111",  "111111011011010110",  "111111011011110100",  "111111011100010011",  "111111011100110001",  "111111011101010000",  "111111011101101111",  "111111011110001101",  "111111011110101100",  "111111011111001010",  "111111011111101001",  "111111100000000111",  "111111100000100110",  "111111100001000101",  "111111100001100011",  "111111100010000010",  "111111100010100000",  "111111100010111111",  "111111100011011110",  "111111100011111100",  "111111100100011011",  "111111100100111001",  "111111100101011000",  "111111100101110111",  "111111100110010101",  "111111100110110100",  "111111100111010010",  "111111100111110001",  "111111101000010000",  "111111101000101110",  "111111101001001101",  "111111101001101011",  "111111101010001010",  "111111101010101001",  "111111101011000111",  "111111101011100110",  "111111101100000100",  "111111101100100011",  "111111101101000001",  "111111101101100000",  "111111101101111110",  "111111101110011101",  "111111101110111011",  "111111101111011010",  "111111101111111001",  "111111110000010111",  "111111110000110110",  "111111110001010100",  "111111110001110011",  "111111110010010001",  "111111110010101111",  "111111110011001110",  "111111110011101100",  "111111110100001011",  "111111110100101001",  "111111110101001000",  "111111110101100110",  "111111110110000100",  "111111110110100011",  "111111110111000001",  "111111110111100000",  "111111110111111110",  "111111111000011100",  "111111111000111011",  "111111111001011001",  "111111111001110111",  "111111111010010110",  "111111111010110100",  "111111111011010010",  "111111111011110000",  "111111111100001111",  "111111111100101101",  "111111111101001011",  "111111111101101001",  "111111111110000111",  "111111111110100110",  "111111111111000100",  "111111111111100010"),("000000000000000000",  "000000000000011110",  "000000000000111100",  "000000000001011010",  "000000000001111000",  "000000000010010110",  "000000000010110100",  "000000000011010010",  "000000000011110000",  "000000000100001110",  "000000000100101100",  "000000000101001010",  "000000000101101000",  "000000000110000110",  "000000000110100100",  "000000000111000010",  "000000000111011111",  "000000000111111101",  "000000001000011011",  "000000001000111001",  "000000001001010111",  "000000001001110100",  "000000001010010010",  "000000001010110000",  "000000001011001101",  "000000001011101011",  "000000001100001000",  "000000001100100110",  "000000001101000100",  "000000001101100001",  "000000001101111111",  "000000001110011100",  "000000001110111010",  "000000001111010111",  "000000001111110100",  "000000010000010010",  "000000010000101111",  "000000010001001101",  "000000010001101010",  "000000010010000111",  "000000010010100100",  "000000010011000010",  "000000010011011111",  "000000010011111100",  "000000010100011001",  "000000010100110110",  "000000010101010011",  "000000010101110000",  "000000010110001101",  "000000010110101010",  "000000010111000111",  "000000010111100100",  "000000011000000001",  "000000011000011110",  "000000011000111011",  "000000011001011000",  "000000011001110100",  "000000011010010001",  "000000011010101110",  "000000011011001011",  "000000011011100111",  "000000011100000100",  "000000011100100001",  "000000011100111101",  "000000011101011010",  "000000011101110110",  "000000011110010011",  "000000011110101111",  "000000011111001011",  "000000011111101000",  "000000100000000100",  "000000100000100000",  "000000100000111101",  "000000100001011001",  "000000100001110101",  "000000100010010001",  "000000100010101101",  "000000100011001001",  "000000100011100101",  "000000100100000001",  "000000100100011101",  "000000100100111001",  "000000100101010101",  "000000100101110001",  "000000100110001101",  "000000100110101001",  "000000100111000100",  "000000100111100000",  "000000100111111100",  "000000101000010111",  "000000101000110011",  "000000101001001111",  "000000101001101010",  "000000101010000101",  "000000101010100001",  "000000101010111100",  "000000101011011000",  "000000101011110011",  "000000101100001110",  "000000101100101001",  "000000101101000101",  "000000101101100000",  "000000101101111011",  "000000101110010110",  "000000101110110001",  "000000101111001100",  "000000101111100111",  "000000110000000010",  "000000110000011101",  "000000110000110111",  "000000110001010010",  "000000110001101101",  "000000110010000111",  "000000110010100010",  "000000110010111101",  "000000110011010111",  "000000110011110010",  "000000110100001100",  "000000110100100110",  "000000110101000001",  "000000110101011011",  "000000110101110101",  "000000110110010000",  "000000110110101010",  "000000110111000100",  "000000110111011110",  "000000110111111000",  "000000111000010010",  "000000111000101100",  "000000111001000110",  "000000111001100000",  "000000111001111001",  "000000111010010011",  "000000111010101101",  "000000111011000110",  "000000111011100000",  "000000111011111001",  "000000111100010011",  "000000111100101100",  "000000111101000110",  "000000111101011111",  "000000111101111000",  "000000111110010010",  "000000111110101011",  "000000111111000100",  "000000111111011101",  "000000111111110110",  "000001000000001111",  "000001000000101000",  "000001000001000001",  "000001000001011010",  "000001000001110010",  "000001000010001011",  "000001000010100100",  "000001000010111100",  "000001000011010101",  "000001000011101101",  "000001000100000110",  "000001000100011110",  "000001000100110111",  "000001000101001111",  "000001000101100111",  "000001000101111111",  "000001000110010111",  "000001000110101111",  "000001000111000111",  "000001000111011111",  "000001000111110111",  "000001001000001111",  "000001001000100111",  "000001001000111111",  "000001001001010110",  "000001001001101110",  "000001001010000101",  "000001001010011101",  "000001001010110100",  "000001001011001100",  "000001001011100011",  "000001001011111010",  "000001001100010010",  "000001001100101001",  "000001001101000000",  "000001001101010111",  "000001001101101110",  "000001001110000101",  "000001001110011100",  "000001001110110010",  "000001001111001001",  "000001001111100000",  "000001001111110110",  "000001010000001101",  "000001010000100011",  "000001010000111010",  "000001010001010000",  "000001010001100111",  "000001010001111101",  "000001010010010011",  "000001010010101001",  "000001010010111111",  "000001010011010101",  "000001010011101011",  "000001010100000001",  "000001010100010111",  "000001010100101101",  "000001010101000010",  "000001010101011000",  "000001010101101110",  "000001010110000011",  "000001010110011000",  "000001010110101110",  "000001010111000011",  "000001010111011000",  "000001010111101110",  "000001011000000011",  "000001011000011000",  "000001011000101101",  "000001011001000010",  "000001011001010111",  "000001011001101011",  "000001011010000000",  "000001011010010101",  "000001011010101001",  "000001011010111110",  "000001011011010010",  "000001011011100111",  "000001011011111011",  "000001011100001111",  "000001011100100100",  "000001011100111000",  "000001011101001100",  "000001011101100000",  "000001011101110100",  "000001011110001000",  "000001011110011011",  "000001011110101111",  "000001011111000011",  "000001011111010111",  "000001011111101010",  "000001011111111110",  "000001100000010001",  "000001100000100100",  "000001100000111000",  "000001100001001011",  "000001100001011110",  "000001100001110001",  "000001100010000100",  "000001100010010111",  "000001100010101010",  "000001100010111100",  "000001100011001111",  "000001100011100010",  "000001100011110100",  "000001100100000111",  "000001100100011001",  "000001100100101100",  "000001100100111110",  "000001100101010000",  "000001100101100010",  "000001100101110100",  "000001100110000110",  "000001100110011000",  "000001100110101010",  "000001100110111100",  "000001100111001110",  "000001100111011111",  "000001100111110001",  "000001101000000010",  "000001101000010100",  "000001101000100101",  "000001101000110111",  "000001101001001000",  "000001101001011001",  "000001101001101010",  "000001101001111011",  "000001101010001100",  "000001101010011101",  "000001101010101110",  "000001101010111110",  "000001101011001111",  "000001101011100000",  "000001101011110000",  "000001101100000000",  "000001101100010001",  "000001101100100001",  "000001101100110001",  "000001101101000001",  "000001101101010001",  "000001101101100001",  "000001101101110001",  "000001101110000001",  "000001101110010001",  "000001101110100000",  "000001101110110000",  "000001101111000000",  "000001101111001111",  "000001101111011110",  "000001101111101110",  "000001101111111101",  "000001110000001100",  "000001110000011011",  "000001110000101010",  "000001110000111001",  "000001110001001000",  "000001110001010111",  "000001110001100101",  "000001110001110100",  "000001110010000011",  "000001110010010001",  "000001110010011111",  "000001110010101110",  "000001110010111100",  "000001110011001010",  "000001110011011000",  "000001110011100110",  "000001110011110100",  "000001110100000010",  "000001110100010000",  "000001110100011101",  "000001110100101011",  "000001110100111001",  "000001110101000110",  "000001110101010011",  "000001110101100001",  "000001110101101110",  "000001110101111011",  "000001110110001000",  "000001110110010101",  "000001110110100010",  "000001110110101111",  "000001110110111100",  "000001110111001000",  "000001110111010101",  "000001110111100010",  "000001110111101110",  "000001110111111010",  "000001111000000111",  "000001111000010011",  "000001111000011111",  "000001111000101011",  "000001111000110111",  "000001111001000011",  "000001111001001111",  "000001111001011010",  "000001111001100110",  "000001111001110010",  "000001111001111101",  "000001111010001001",  "000001111010010100",  "000001111010011111",  "000001111010101010",  "000001111010110101",  "000001111011000000",  "000001111011001011",  "000001111011010110",  "000001111011100001",  "000001111011101100",  "000001111011110110",  "000001111100000001",  "000001111100001011",  "000001111100010110",  "000001111100100000",  "000001111100101010",  "000001111100110100",  "000001111100111110",  "000001111101001000",  "000001111101010010",  "000001111101011100",  "000001111101100110",  "000001111101110000",  "000001111101111001",  "000001111110000011",  "000001111110001100",  "000001111110010101",  "000001111110011111",  "000001111110101000",  "000001111110110001",  "000001111110111010",  "000001111111000011",  "000001111111001100",  "000001111111010100",  "000001111111011101",  "000001111111100110",  "000001111111101110",  "000001111111110111",  "000001111111111111",  "000010000000000111",  "000010000000001111",  "000010000000010111",  "000010000000100000",  "000010000000100111",  "000010000000101111",  "000010000000110111",  "000010000000111111",  "000010000001000110",  "000010000001001110",  "000010000001010101",  "000010000001011101",  "000010000001100100",  "000010000001101011",  "000010000001110010",  "000010000001111001",  "000010000010000000",  "000010000010000111",  "000010000010001110",  "000010000010010101",  "000010000010011011",  "000010000010100010",  "000010000010101000",  "000010000010101111",  "000010000010110101",  "000010000010111011",  "000010000011000010",  "000010000011001000",  "000010000011001110",  "000010000011010011",  "000010000011011001",  "000010000011011111",  "000010000011100101",  "000010000011101010",  "000010000011110000",  "000010000011110101",  "000010000011111010",  "000010000100000000",  "000010000100000101",  "000010000100001010",  "000010000100001111",  "000010000100010100",  "000010000100011001",  "000010000100011101",  "000010000100100010",  "000010000100100111",  "000010000100101011",  "000010000100101111",  "000010000100110100",  "000010000100111000",  "000010000100111100",  "000010000101000000",  "000010000101000100",  "000010000101001000",  "000010000101001100",  "000010000101010000",  "000010000101010011",  "000010000101010111",  "000010000101011011",  "000010000101011110",  "000010000101100001",  "000010000101100101",  "000010000101101000",  "000010000101101011",  "000010000101101110",  "000010000101110001",  "000010000101110100",  "000010000101110110",  "000010000101111001",  "000010000101111100",  "000010000101111110",  "000010000110000001",  "000010000110000011",  "000010000110000101",  "000010000110000111",  "000010000110001010",  "000010000110001100",  "000010000110001110",  "000010000110001111",  "000010000110010001",  "000010000110010011",  "000010000110010101",  "000010000110010110",  "000010000110011000",  "000010000110011001",  "000010000110011010",  "000010000110011011",  "000010000110011101",  "000010000110011110",  "000010000110011111",  "000010000110011111",  "000010000110100000",  "000010000110100001",  "000010000110100010",  "000010000110100010",  "000010000110100011",  "000010000110100011",  "000010000110100011",  "000010000110100011",  "000010000110100100",  "000010000110100100",  "000010000110100100",  "000010000110100100",  "000010000110100011",  "000010000110100011",  "000010000110100011",  "000010000110100010",  "000010000110100010",  "000010000110100001",  "000010000110100001",  "000010000110100000",  "000010000110011111",  "000010000110011110",  "000010000110011101",  "000010000110011100",  "000010000110011011",  "000010000110011010",  "000010000110011000",  "000010000110010111",  "000010000110010110",  "000010000110010100",  "000010000110010010",  "000010000110010001",  "000010000110001111",  "000010000110001101",  "000010000110001011",  "000010000110001001",  "000010000110000111",  "000010000110000101",  "000010000110000010",  "000010000110000000",  "000010000101111110",  "000010000101111011",  "000010000101111001",  "000010000101110110",  "000010000101110011",  "000010000101110000",  "000010000101101101",  "000010000101101010",  "000010000101100111",  "000010000101100100",  "000010000101100001",  "000010000101011110",  "000010000101011010",  "000010000101010111",  "000010000101010011",  "000010000101010000",  "000010000101001100",  "000010000101001000",  "000010000101000100",  "000010000101000000",  "000010000100111100",  "000010000100111000",  "000010000100110100",  "000010000100110000",  "000010000100101100",  "000010000100100111",  "000010000100100011",  "000010000100011110",  "000010000100011001",  "000010000100010101",  "000010000100010000",  "000010000100001011",  "000010000100000110",  "000010000100000001",  "000010000011111100",  "000010000011110111",  "000010000011110010",  "000010000011101100",  "000010000011100111",  "000010000011100001",  "000010000011011100",  "000010000011010110",  "000010000011010000",  "000010000011001011",  "000010000011000101",  "000010000010111111",  "000010000010111001",  "000010000010110011",  "000010000010101101",  "000010000010100110",  "000010000010100000",  "000010000010011010",  "000010000010010011",  "000010000010001101",  "000010000010000110",  "000010000001111111",  "000010000001111000",  "000010000001110010",  "000010000001101011",  "000010000001100100",  "000010000001011101",  "000010000001010101",  "000010000001001110",  "000010000001000111",  "000010000001000000",  "000010000000111000",  "000010000000110001",  "000010000000101001",  "000010000000100001",  "000010000000011010",  "000010000000010010",  "000010000000001010",  "000010000000000010",  "000001111111111010",  "000001111111110010",  "000001111111101010",  "000001111111100001",  "000001111111011001",  "000001111111010001",  "000001111111001000",  "000001111111000000",  "000001111110110111",  "000001111110101110",  "000001111110100110",  "000001111110011101",  "000001111110010100",  "000001111110001011",  "000001111110000010",  "000001111101111001",  "000001111101101111",  "000001111101100110",  "000001111101011101",  "000001111101010011",  "000001111101001010",  "000001111101000000",  "000001111100110111",  "000001111100101101",  "000001111100100011",  "000001111100011001",  "000001111100010000",  "000001111100000110",  "000001111011111100",  "000001111011110001",  "000001111011100111",  "000001111011011101",  "000001111011010011",  "000001111011001000",  "000001111010111110",  "000001111010110011",  "000001111010101001",  "000001111010011110",  "000001111010010011",  "000001111010001000",  "000001111001111110",  "000001111001110011",  "000001111001101000",  "000001111001011101",  "000001111001010001",  "000001111001000110",  "000001111000111011",  "000001111000110000",  "000001111000100100",  "000001111000011001",  "000001111000001101",  "000001111000000010",  "000001110111110110",  "000001110111101010",  "000001110111011110",  "000001110111010010",  "000001110111000110",  "000001110110111010",  "000001110110101110",  "000001110110100010",  "000001110110010110",  "000001110110001010",  "000001110101111101",  "000001110101110001",  "000001110101100100",  "000001110101011000",  "000001110101001011",  "000001110100111111",  "000001110100110010",  "000001110100100101",  "000001110100011000",  "000001110100001011",  "000001110011111110",  "000001110011110001",  "000001110011100100",  "000001110011010111",  "000001110011001010",  "000001110010111100",  "000001110010101111",  "000001110010100010",  "000001110010010100",  "000001110010000111",  "000001110001111001",  "000001110001101011",  "000001110001011110",  "000001110001010000",  "000001110001000010",  "000001110000110100",  "000001110000100110",  "000001110000011000",  "000001110000001010",  "000001101111111100",  "000001101111101101",  "000001101111011111",  "000001101111010001",  "000001101111000010",  "000001101110110100",  "000001101110100101",  "000001101110010111",  "000001101110001000",  "000001101101111001",  "000001101101101011",  "000001101101011100",  "000001101101001101",  "000001101100111110",  "000001101100101111",  "000001101100100000",  "000001101100010001",  "000001101100000010",  "000001101011110010",  "000001101011100011",  "000001101011010100",  "000001101011000100",  "000001101010110101",  "000001101010100101",  "000001101010010110",  "000001101010000110",  "000001101001110110",  "000001101001100111",  "000001101001010111",  "000001101001000111",  "000001101000110111",  "000001101000100111",  "000001101000010111",  "000001101000000111",  "000001100111110111",  "000001100111100111",  "000001100111010110",  "000001100111000110",  "000001100110110110",  "000001100110100101",  "000001100110010101",  "000001100110000100",  "000001100101110100",  "000001100101100011",  "000001100101010011",  "000001100101000010",  "000001100100110001",  "000001100100100000",  "000001100100001111",  "000001100011111110",  "000001100011101101",  "000001100011011100",  "000001100011001011",  "000001100010111010",  "000001100010101001",  "000001100010011000",  "000001100010000110",  "000001100001110101",  "000001100001100100",  "000001100001010010",  "000001100001000001",  "000001100000101111",  "000001100000011101",  "000001100000001100",  "000001011111111010",  "000001011111101000",  "000001011111010110",  "000001011111000101",  "000001011110110011",  "000001011110100001",  "000001011110001111",  "000001011101111101",  "000001011101101011",  "000001011101011000",  "000001011101000110",  "000001011100110100",  "000001011100100010",  "000001011100001111",  "000001011011111101",  "000001011011101011",  "000001011011011000",  "000001011011000110",  "000001011010110011",  "000001011010100000",  "000001011010001110",  "000001011001111011",  "000001011001101000",  "000001011001010110",  "000001011001000011",  "000001011000110000",  "000001011000011101",  "000001011000001010",  "000001010111110111",  "000001010111100100",  "000001010111010001",  "000001010110111110",  "000001010110101010",  "000001010110010111",  "000001010110000100",  "000001010101110001",  "000001010101011101",  "000001010101001010",  "000001010100110110",  "000001010100100011",  "000001010100001111",  "000001010011111100",  "000001010011101000",  "000001010011010101",  "000001010011000001",  "000001010010101101",  "000001010010011001",  "000001010010000110",  "000001010001110010",  "000001010001011110",  "000001010001001010",  "000001010000110110",  "000001010000100010",  "000001010000001110",  "000001001111111010",  "000001001111100110",  "000001001111010010",  "000001001110111101",  "000001001110101001",  "000001001110010101",  "000001001110000000",  "000001001101101100",  "000001001101011000",  "000001001101000011",  "000001001100101111",  "000001001100011010",  "000001001100000110",  "000001001011110001",  "000001001011011101",  "000001001011001000",  "000001001010110011",  "000001001010011111",  "000001001010001010",  "000001001001110101",  "000001001001100000",  "000001001001001011",  "000001001000110110",  "000001001000100010",  "000001001000001101",  "000001000111111000",  "000001000111100011",  "000001000111001101",  "000001000110111000",  "000001000110100011",  "000001000110001110",  "000001000101111001",  "000001000101100100",  "000001000101001110",  "000001000100111001",  "000001000100100100",  "000001000100001111",  "000001000011111001",  "000001000011100100",  "000001000011001110",  "000001000010111001",  "000001000010100011",  "000001000010001110",  "000001000001111000",  "000001000001100011",  "000001000001001101",  "000001000000110111",  "000001000000100010",  "000001000000001100",  "000000111111110110",  "000000111111100001",  "000000111111001011",  "000000111110110101",  "000000111110011111",  "000000111110001001",  "000000111101110011",  "000000111101011101",  "000000111101000111",  "000000111100110001",  "000000111100011011",  "000000111100000101",  "000000111011101111",  "000000111011011001",  "000000111011000011",  "000000111010101101",  "000000111010010111",  "000000111010000001",  "000000111001101011",  "000000111001010100",  "000000111000111110",  "000000111000101000",  "000000111000010001",  "000000110111111011",  "000000110111100101",  "000000110111001110",  "000000110110111000",  "000000110110100010",  "000000110110001011",  "000000110101110101",  "000000110101011110",  "000000110101001000",  "000000110100110001",  "000000110100011011",  "000000110100000100",  "000000110011101101",  "000000110011010111",  "000000110011000000",  "000000110010101010",  "000000110010010011",  "000000110001111100",  "000000110001100110",  "000000110001001111",  "000000110000111000",  "000000110000100001",  "000000110000001010",  "000000101111110100",  "000000101111011101",  "000000101111000110",  "000000101110101111",  "000000101110011000",  "000000101110000001",  "000000101101101011",  "000000101101010100",  "000000101100111101",  "000000101100100110",  "000000101100001111",  "000000101011111000",  "000000101011100001",  "000000101011001010",  "000000101010110011",  "000000101010011100",  "000000101010000101",  "000000101001101101",  "000000101001010110",  "000000101000111111",  "000000101000101000",  "000000101000010001",  "000000100111111010",  "000000100111100011",  "000000100111001100",  "000000100110110100",  "000000100110011101",  "000000100110000110",  "000000100101101111",  "000000100101011000",  "000000100101000000",  "000000100100101001",  "000000100100010010",  "000000100011111010",  "000000100011100011",  "000000100011001100",  "000000100010110101",  "000000100010011101",  "000000100010000110",  "000000100001101111",  "000000100001010111",  "000000100001000000",  "000000100000101000",  "000000100000010001",  "000000011111111010",  "000000011111100010",  "000000011111001011",  "000000011110110100",  "000000011110011100",  "000000011110000101",  "000000011101101101",  "000000011101010110",  "000000011100111110",  "000000011100100111",  "000000011100001111",  "000000011011111000",  "000000011011100001",  "000000011011001001",  "000000011010110010",  "000000011010011010",  "000000011010000011",  "000000011001101011",  "000000011001010100",  "000000011000111100",  "000000011000100101",  "000000011000001101",  "000000010111110110",  "000000010111011110",  "000000010111000111",  "000000010110101111",  "000000010110010111",  "000000010110000000",  "000000010101101000",  "000000010101010001",  "000000010100111001",  "000000010100100010",  "000000010100001010",  "000000010011110011",  "000000010011011011",  "000000010011000100",  "000000010010101100",  "000000010010010101",  "000000010001111101",  "000000010001100101",  "000000010001001110",  "000000010000110110",  "000000010000011111",  "000000010000000111",  "000000001111110000",  "000000001111011000",  "000000001111000001",  "000000001110101001",  "000000001110010010",  "000000001101111010",  "000000001101100011",  "000000001101001011",  "000000001100110100",  "000000001100011100",  "000000001100000101",  "000000001011101101",  "000000001011010110",  "000000001010111110",  "000000001010100111",  "000000001010001111",  "000000001001111000",  "000000001001100000",  "000000001001001001",  "000000001000110001",  "000000001000011010",  "000000001000000010",  "000000000111101011",  "000000000111010011",  "000000000110111100",  "000000000110100100",  "000000000110001101",  "000000000101110110",  "000000000101011110",  "000000000101000111",  "000000000100101111",  "000000000100011000",  "000000000100000001",  "000000000011101001",  "000000000011010010",  "000000000010111010",  "000000000010100011",  "000000000010001100",  "000000000001110100",  "000000000001011101",  "000000000001000110",  "000000000000101111",  "000000000000010111"),("000000000000000000",  "111111111111101001",  "111111111111010001",  "111111111110111010",  "111111111110100011",  "111111111110001100",  "111111111101110101",  "111111111101011101",  "111111111101000110",  "111111111100101111",  "111111111100011000",  "111111111100000001",  "111111111011101010",  "111111111011010010",  "111111111010111011",  "111111111010100100",  "111111111010001101",  "111111111001110110",  "111111111001011111",  "111111111001001000",  "111111111000110001",  "111111111000011010",  "111111111000000011",  "111111110111101100",  "111111110111010101",  "111111110110111110",  "111111110110100111",  "111111110110010000",  "111111110101111001",  "111111110101100011",  "111111110101001100",  "111111110100110101",  "111111110100011110",  "111111110100000111",  "111111110011110000",  "111111110011011010",  "111111110011000011",  "111111110010101100",  "111111110010010110",  "111111110001111111",  "111111110001101000",  "111111110001010001",  "111111110000111011",  "111111110000100100",  "111111110000001110",  "111111101111110111",  "111111101111100000",  "111111101111001010",  "111111101110110011",  "111111101110011101",  "111111101110000110",  "111111101101110000",  "111111101101011010",  "111111101101000011",  "111111101100101101",  "111111101100010110",  "111111101100000000",  "111111101011101010",  "111111101011010011",  "111111101010111101",  "111111101010100111",  "111111101010010001",  "111111101001111010",  "111111101001100100",  "111111101001001110",  "111111101000111000",  "111111101000100010",  "111111101000001100",  "111111100111110110",  "111111100111100000",  "111111100111001010",  "111111100110110100",  "111111100110011110",  "111111100110001000",  "111111100101110010",  "111111100101011100",  "111111100101000110",  "111111100100110000",  "111111100100011010",  "111111100100000101",  "111111100011101111",  "111111100011011001",  "111111100011000011",  "111111100010101110",  "111111100010011000",  "111111100010000011",  "111111100001101101",  "111111100001010111",  "111111100001000010",  "111111100000101100",  "111111100000010111",  "111111100000000001",  "111111011111101100",  "111111011111010111",  "111111011111000001",  "111111011110101100",  "111111011110010111",  "111111011110000001",  "111111011101101100",  "111111011101010111",  "111111011101000010",  "111111011100101101",  "111111011100010111",  "111111011100000010",  "111111011011101101",  "111111011011011000",  "111111011011000011",  "111111011010101110",  "111111011010011001",  "111111011010000101",  "111111011001110000",  "111111011001011011",  "111111011001000110",  "111111011000110001",  "111111011000011101",  "111111011000001000",  "111111010111110011",  "111111010111011111",  "111111010111001010",  "111111010110110101",  "111111010110100001",  "111111010110001100",  "111111010101111000",  "111111010101100100",  "111111010101001111",  "111111010100111011",  "111111010100100111",  "111111010100010010",  "111111010011111110",  "111111010011101010",  "111111010011010110",  "111111010011000001",  "111111010010101101",  "111111010010011001",  "111111010010000101",  "111111010001110001",  "111111010001011101",  "111111010001001001",  "111111010000110110",  "111111010000100010",  "111111010000001110",  "111111001111111010",  "111111001111100110",  "111111001111010011",  "111111001110111111",  "111111001110101011",  "111111001110011000",  "111111001110000100",  "111111001101110001",  "111111001101011101",  "111111001101001010",  "111111001100110111",  "111111001100100011",  "111111001100010000",  "111111001011111101",  "111111001011101010",  "111111001011010110",  "111111001011000011",  "111111001010110000",  "111111001010011101",  "111111001010001010",  "111111001001110111",  "111111001001100100",  "111111001001010001",  "111111001000111110",  "111111001000101100",  "111111001000011001",  "111111001000000110",  "111111000111110011",  "111111000111100001",  "111111000111001110",  "111111000110111100",  "111111000110101001",  "111111000110010111",  "111111000110000100",  "111111000101110010",  "111111000101100000",  "111111000101001101",  "111111000100111011",  "111111000100101001",  "111111000100010111",  "111111000100000101",  "111111000011110010",  "111111000011100000",  "111111000011001110",  "111111000010111100",  "111111000010101011",  "111111000010011001",  "111111000010000111",  "111111000001110101",  "111111000001100011",  "111111000001010010",  "111111000001000000",  "111111000000101111",  "111111000000011101",  "111111000000001100",  "111110111111111010",  "111110111111101001",  "111110111111010111",  "111110111111000110",  "111110111110110101",  "111110111110100100",  "111110111110010011",  "111110111110000001",  "111110111101110000",  "111110111101011111",  "111110111101001110",  "111110111100111110",  "111110111100101101",  "111110111100011100",  "111110111100001011",  "111110111011111010",  "111110111011101010",  "111110111011011001",  "111110111011001000",  "111110111010111000",  "111110111010101000",  "111110111010010111",  "111110111010000111",  "111110111001110110",  "111110111001100110",  "111110111001010110",  "111110111001000110",  "111110111000110110",  "111110111000100101",  "111110111000010101",  "111110111000000101",  "111110110111110110",  "111110110111100110",  "111110110111010110",  "111110110111000110",  "111110110110110110",  "111110110110100111",  "111110110110010111",  "111110110110001000",  "111110110101111000",  "111110110101101001",  "111110110101011001",  "111110110101001010",  "111110110100111010",  "111110110100101011",  "111110110100011100",  "111110110100001101",  "111110110011111110",  "111110110011101111",  "111110110011100000",  "111110110011010001",  "111110110011000010",  "111110110010110011",  "111110110010100100",  "111110110010010110",  "111110110010000111",  "111110110001111000",  "111110110001101010",  "111110110001011011",  "111110110001001101",  "111110110000111110",  "111110110000110000",  "111110110000100010",  "111110110000010011",  "111110110000000101",  "111110101111110111",  "111110101111101001",  "111110101111011011",  "111110101111001101",  "111110101110111111",  "111110101110110001",  "111110101110100100",  "111110101110010110",  "111110101110001000",  "111110101101111010",  "111110101101101101",  "111110101101011111",  "111110101101010010",  "111110101101000100",  "111110101100110111",  "111110101100101010",  "111110101100011101",  "111110101100001111",  "111110101100000010",  "111110101011110101",  "111110101011101000",  "111110101011011011",  "111110101011001110",  "111110101011000001",  "111110101010110101",  "111110101010101000",  "111110101010011011",  "111110101010001111",  "111110101010000010",  "111110101001110110",  "111110101001101001",  "111110101001011101",  "111110101001010000",  "111110101001000100",  "111110101000111000",  "111110101000101100",  "111110101000100000",  "111110101000010100",  "111110101000001000",  "111110100111111100",  "111110100111110000",  "111110100111100100",  "111110100111011000",  "111110100111001101",  "111110100111000001",  "111110100110110101",  "111110100110101010",  "111110100110011110",  "111110100110010011",  "111110100110001000",  "111110100101111101",  "111110100101110001",  "111110100101100110",  "111110100101011011",  "111110100101010000",  "111110100101000101",  "111110100100111010",  "111110100100101111",  "111110100100100100",  "111110100100011010",  "111110100100001111",  "111110100100000100",  "111110100011111010",  "111110100011101111",  "111110100011100101",  "111110100011011011",  "111110100011010000",  "111110100011000110",  "111110100010111100",  "111110100010110010",  "111110100010101000",  "111110100010011110",  "111110100010010100",  "111110100010001010",  "111110100010000000",  "111110100001110110",  "111110100001101100",  "111110100001100011",  "111110100001011001",  "111110100001010000",  "111110100001000110",  "111110100000111101",  "111110100000110100",  "111110100000101010",  "111110100000100001",  "111110100000011000",  "111110100000001111",  "111110100000000110",  "111110011111111101",  "111110011111110100",  "111110011111101011",  "111110011111100010",  "111110011111011010",  "111110011111010001",  "111110011111001000",  "111110011111000000",  "111110011110110111",  "111110011110101111",  "111110011110100111",  "111110011110011110",  "111110011110010110",  "111110011110001110",  "111110011110000110",  "111110011101111110",  "111110011101110110",  "111110011101101110",  "111110011101100110",  "111110011101011110",  "111110011101010111",  "111110011101001111",  "111110011101000111",  "111110011101000000",  "111110011100111000",  "111110011100110001",  "111110011100101010",  "111110011100100010",  "111110011100011011",  "111110011100010100",  "111110011100001101",  "111110011100000110",  "111110011011111111",  "111110011011111000",  "111110011011110001",  "111110011011101011",  "111110011011100100",  "111110011011011101",  "111110011011010111",  "111110011011010000",  "111110011011001010",  "111110011011000011",  "111110011010111101",  "111110011010110111",  "111110011010110001",  "111110011010101010",  "111110011010100100",  "111110011010011110",  "111110011010011000",  "111110011010010011",  "111110011010001101",  "111110011010000111",  "111110011010000001",  "111110011001111100",  "111110011001110110",  "111110011001110001",  "111110011001101011",  "111110011001100110",  "111110011001100001",  "111110011001011011",  "111110011001010110",  "111110011001010001",  "111110011001001100",  "111110011001000111",  "111110011001000010",  "111110011000111101",  "111110011000111000",  "111110011000110100",  "111110011000101111",  "111110011000101011",  "111110011000100110",  "111110011000100010",  "111110011000011101",  "111110011000011001",  "111110011000010101",  "111110011000010000",  "111110011000001100",  "111110011000001000",  "111110011000000100",  "111110011000000000",  "111110010111111100",  "111110010111111001",  "111110010111110101",  "111110010111110001",  "111110010111101101",  "111110010111101010",  "111110010111100110",  "111110010111100011",  "111110010111100000",  "111110010111011100",  "111110010111011001",  "111110010111010110",  "111110010111010011",  "111110010111010000",  "111110010111001101",  "111110010111001010",  "111110010111000111",  "111110010111000100",  "111110010111000010",  "111110010110111111",  "111110010110111100",  "111110010110111010",  "111110010110110111",  "111110010110110101",  "111110010110110011",  "111110010110110000",  "111110010110101110",  "111110010110101100",  "111110010110101010",  "111110010110101000",  "111110010110100110",  "111110010110100100",  "111110010110100010",  "111110010110100001",  "111110010110011111",  "111110010110011101",  "111110010110011100",  "111110010110011010",  "111110010110011001",  "111110010110010111",  "111110010110010110",  "111110010110010101",  "111110010110010100",  "111110010110010011",  "111110010110010010",  "111110010110010001",  "111110010110010000",  "111110010110001111",  "111110010110001110",  "111110010110001101",  "111110010110001101",  "111110010110001100",  "111110010110001100",  "111110010110001011",  "111110010110001011",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001010",  "111110010110001011",  "111110010110001011",  "111110010110001011",  "111110010110001100",  "111110010110001100",  "111110010110001101",  "111110010110001110",  "111110010110001111",  "111110010110001111",  "111110010110010000",  "111110010110010001",  "111110010110010010",  "111110010110010011",  "111110010110010100",  "111110010110010110",  "111110010110010111",  "111110010110011000",  "111110010110011010",  "111110010110011011",  "111110010110011101",  "111110010110011110",  "111110010110100000",  "111110010110100001",  "111110010110100011",  "111110010110100101",  "111110010110100111",  "111110010110101001",  "111110010110101011",  "111110010110101101",  "111110010110101111",  "111110010110110001",  "111110010110110100",  "111110010110110110",  "111110010110111000",  "111110010110111011",  "111110010110111101",  "111110010111000000",  "111110010111000010",  "111110010111000101",  "111110010111001000",  "111110010111001011",  "111110010111001110",  "111110010111010001",  "111110010111010100",  "111110010111010111",  "111110010111011010",  "111110010111011101",  "111110010111100000",  "111110010111100100",  "111110010111100111",  "111110010111101010",  "111110010111101110",  "111110010111110001",  "111110010111110101",  "111110010111111001",  "111110010111111101",  "111110011000000000",  "111110011000000100",  "111110011000001000",  "111110011000001100",  "111110011000010000",  "111110011000010100",  "111110011000011001",  "111110011000011101",  "111110011000100001",  "111110011000100101",  "111110011000101010",  "111110011000101110",  "111110011000110011",  "111110011000110111",  "111110011000111100",  "111110011001000001",  "111110011001000110",  "111110011001001010",  "111110011001001111",  "111110011001010100",  "111110011001011001",  "111110011001011110",  "111110011001100100",  "111110011001101001",  "111110011001101110",  "111110011001110011",  "111110011001111001",  "111110011001111110",  "111110011010000100",  "111110011010001001",  "111110011010001111",  "111110011010010101",  "111110011010011010",  "111110011010100000",  "111110011010100110",  "111110011010101100",  "111110011010110010",  "111110011010111000",  "111110011010111110",  "111110011011000100",  "111110011011001010",  "111110011011010001",  "111110011011010111",  "111110011011011101",  "111110011011100100",  "111110011011101010",  "111110011011110001",  "111110011011110111",  "111110011011111110",  "111110011100000101",  "111110011100001100",  "111110011100010010",  "111110011100011001",  "111110011100100000",  "111110011100100111",  "111110011100101110",  "111110011100110101",  "111110011100111101",  "111110011101000100",  "111110011101001011",  "111110011101010010",  "111110011101011010",  "111110011101100001",  "111110011101101001",  "111110011101110000",  "111110011101111000",  "111110011110000000",  "111110011110001000",  "111110011110001111",  "111110011110010111",  "111110011110011111",  "111110011110100111",  "111110011110101111",  "111110011110110111",  "111110011110111111",  "111110011111000111",  "111110011111010000",  "111110011111011000",  "111110011111100000",  "111110011111101001",  "111110011111110001",  "111110011111111010",  "111110100000000010",  "111110100000001011",  "111110100000010100",  "111110100000011100",  "111110100000100101",  "111110100000101110",  "111110100000110111",  "111110100001000000",  "111110100001001001",  "111110100001010010",  "111110100001011011",  "111110100001100100",  "111110100001101101",  "111110100001110111",  "111110100010000000",  "111110100010001001",  "111110100010010011",  "111110100010011100",  "111110100010100110",  "111110100010101111",  "111110100010111001",  "111110100011000011",  "111110100011001100",  "111110100011010110",  "111110100011100000",  "111110100011101010",  "111110100011110100",  "111110100011111110",  "111110100100001000",  "111110100100010010",  "111110100100011100",  "111110100100100110",  "111110100100110001",  "111110100100111011",  "111110100101000101",  "111110100101010000",  "111110100101011010",  "111110100101100101",  "111110100101101111",  "111110100101111010",  "111110100110000100",  "111110100110001111",  "111110100110011010",  "111110100110100101",  "111110100110110000",  "111110100110111010",  "111110100111000101",  "111110100111010000",  "111110100111011011",  "111110100111100110",  "111110100111110010",  "111110100111111101",  "111110101000001000",  "111110101000010011",  "111110101000011111",  "111110101000101010",  "111110101000110110",  "111110101001000001",  "111110101001001101",  "111110101001011000",  "111110101001100100",  "111110101001101111",  "111110101001111011",  "111110101010000111",  "111110101010010011",  "111110101010011111",  "111110101010101010",  "111110101010110110",  "111110101011000010",  "111110101011001110",  "111110101011011011",  "111110101011100111",  "111110101011110011",  "111110101011111111",  "111110101100001011",  "111110101100011000",  "111110101100100100",  "111110101100110000",  "111110101100111101",  "111110101101001001",  "111110101101010110",  "111110101101100011",  "111110101101101111",  "111110101101111100",  "111110101110001001",  "111110101110010101",  "111110101110100010",  "111110101110101111",  "111110101110111100",  "111110101111001001",  "111110101111010110",  "111110101111100011",  "111110101111110000",  "111110101111111101",  "111110110000001010",  "111110110000010111",  "111110110000100101",  "111110110000110010",  "111110110000111111",  "111110110001001101",  "111110110001011010",  "111110110001100111",  "111110110001110101",  "111110110010000010",  "111110110010010000",  "111110110010011110",  "111110110010101011",  "111110110010111001",  "111110110011000111",  "111110110011010100",  "111110110011100010",  "111110110011110000",  "111110110011111110",  "111110110100001100",  "111110110100011010",  "111110110100101000",  "111110110100110110",  "111110110101000100",  "111110110101010010",  "111110110101100000",  "111110110101101111",  "111110110101111101",  "111110110110001011",  "111110110110011010",  "111110110110101000",  "111110110110110110",  "111110110111000101",  "111110110111010011",  "111110110111100010",  "111110110111110000",  "111110110111111111",  "111110111000001110",  "111110111000011100",  "111110111000101011",  "111110111000111010",  "111110111001001000",  "111110111001010111",  "111110111001100110",  "111110111001110101",  "111110111010000100",  "111110111010010011",  "111110111010100010",  "111110111010110001",  "111110111011000000",  "111110111011001111",  "111110111011011110",  "111110111011101101",  "111110111011111101",  "111110111100001100",  "111110111100011011",  "111110111100101010",  "111110111100111010",  "111110111101001001",  "111110111101011001",  "111110111101101000",  "111110111101110111",  "111110111110000111",  "111110111110010111",  "111110111110100110",  "111110111110110110",  "111110111111000101",  "111110111111010101",  "111110111111100101",  "111110111111110101",  "111111000000000100",  "111111000000010100",  "111111000000100100",  "111111000000110100",  "111111000001000100",  "111111000001010100",  "111111000001100100",  "111111000001110100",  "111111000010000100",  "111111000010010100",  "111111000010100100",  "111111000010110100",  "111111000011000100",  "111111000011010100",  "111111000011100100",  "111111000011110101",  "111111000100000101",  "111111000100010101",  "111111000100100101",  "111111000100110110",  "111111000101000110",  "111111000101010111",  "111111000101100111",  "111111000101111000",  "111111000110001000",  "111111000110011001",  "111111000110101001",  "111111000110111010",  "111111000111001010",  "111111000111011011",  "111111000111101100",  "111111000111111100",  "111111001000001101",  "111111001000011110",  "111111001000101110",  "111111001000111111",  "111111001001010000",  "111111001001100001",  "111111001001110010",  "111111001010000011",  "111111001010010100",  "111111001010100101",  "111111001010110110",  "111111001011000111",  "111111001011011000",  "111111001011101001",  "111111001011111010",  "111111001100001011",  "111111001100011100",  "111111001100101101",  "111111001100111110",  "111111001101001111",  "111111001101100001",  "111111001101110010",  "111111001110000011",  "111111001110010100",  "111111001110100110",  "111111001110110111",  "111111001111001000",  "111111001111011010",  "111111001111101011",  "111111001111111101",  "111111010000001110",  "111111010000011111",  "111111010000110001",  "111111010001000010",  "111111010001010100",  "111111010001100101",  "111111010001110111",  "111111010010001001",  "111111010010011010",  "111111010010101100",  "111111010010111101",  "111111010011001111",  "111111010011100001",  "111111010011110011",  "111111010100000100",  "111111010100010110",  "111111010100101000",  "111111010100111010",  "111111010101001011",  "111111010101011101",  "111111010101101111",  "111111010110000001",  "111111010110010011",  "111111010110100101",  "111111010110110110",  "111111010111001000",  "111111010111011010",  "111111010111101100",  "111111010111111110",  "111111011000010000",  "111111011000100010",  "111111011000110100",  "111111011001000110",  "111111011001011000",  "111111011001101010",  "111111011001111101",  "111111011010001111",  "111111011010100001",  "111111011010110011",  "111111011011000101",  "111111011011010111",  "111111011011101001",  "111111011011111100",  "111111011100001110",  "111111011100100000",  "111111011100110010",  "111111011101000100",  "111111011101010111",  "111111011101101001",  "111111011101111011",  "111111011110001110",  "111111011110100000",  "111111011110110010",  "111111011111000101",  "111111011111010111",  "111111011111101001",  "111111011111111100",  "111111100000001110",  "111111100000100000",  "111111100000110011",  "111111100001000101",  "111111100001011000",  "111111100001101010",  "111111100001111101",  "111111100010001111",  "111111100010100001",  "111111100010110100",  "111111100011000110",  "111111100011011001",  "111111100011101011",  "111111100011111110",  "111111100100010000",  "111111100100100011",  "111111100100110110",  "111111100101001000",  "111111100101011011",  "111111100101101101",  "111111100110000000",  "111111100110010010",  "111111100110100101",  "111111100110111000",  "111111100111001010",  "111111100111011101",  "111111100111101111",  "111111101000000010",  "111111101000010101",  "111111101000100111",  "111111101000111010",  "111111101001001101",  "111111101001011111",  "111111101001110010",  "111111101010000101",  "111111101010010111",  "111111101010101010",  "111111101010111101",  "111111101011001111",  "111111101011100010",  "111111101011110101",  "111111101100000111",  "111111101100011010",  "111111101100101101",  "111111101101000000",  "111111101101010010",  "111111101101100101",  "111111101101111000",  "111111101110001011",  "111111101110011101",  "111111101110110000",  "111111101111000011",  "111111101111010101",  "111111101111101000",  "111111101111111011",  "111111110000001110",  "111111110000100000",  "111111110000110011",  "111111110001000110",  "111111110001011001",  "111111110001101011",  "111111110001111110",  "111111110010010001",  "111111110010100100",  "111111110010110110",  "111111110011001001",  "111111110011011100",  "111111110011101111",  "111111110100000010",  "111111110100010100",  "111111110100100111",  "111111110100111010",  "111111110101001101",  "111111110101011111",  "111111110101110010",  "111111110110000101",  "111111110110011000",  "111111110110101010",  "111111110110111101",  "111111110111010000",  "111111110111100011",  "111111110111110101",  "111111111000001000",  "111111111000011011",  "111111111000101101",  "111111111001000000",  "111111111001010011",  "111111111001100110",  "111111111001111000",  "111111111010001011",  "111111111010011110",  "111111111010110000",  "111111111011000011",  "111111111011010110",  "111111111011101000",  "111111111011111011",  "111111111100001110",  "111111111100100000",  "111111111100110011",  "111111111101000110",  "111111111101011000",  "111111111101101011",  "111111111101111110",  "111111111110010000",  "111111111110100011",  "111111111110110110",  "111111111111001000",  "111111111111011011",  "111111111111101101"),("000000000000000000",  "000000000000010011",  "000000000000100101",  "000000000000111000",  "000000000001001010",  "000000000001011101",  "000000000001101111",  "000000000010000010",  "000000000010010100",  "000000000010100111",  "000000000010111001",  "000000000011001100",  "000000000011011110",  "000000000011110001",  "000000000100000011",  "000000000100010110",  "000000000100101000",  "000000000100111011",  "000000000101001101",  "000000000101100000",  "000000000101110010",  "000000000110000100",  "000000000110010111",  "000000000110101001",  "000000000110111011",  "000000000111001110",  "000000000111100000",  "000000000111110010",  "000000001000000101",  "000000001000010111",  "000000001000101001",  "000000001000111100",  "000000001001001110",  "000000001001100000",  "000000001001110010",  "000000001010000100",  "000000001010010111",  "000000001010101001",  "000000001010111011",  "000000001011001101",  "000000001011011111",  "000000001011110001",  "000000001100000100",  "000000001100010110",  "000000001100101000",  "000000001100111010",  "000000001101001100",  "000000001101011110",  "000000001101110000",  "000000001110000010",  "000000001110010100",  "000000001110100110",  "000000001110111000",  "000000001111001010",  "000000001111011100",  "000000001111101110",  "000000010000000000",  "000000010000010010",  "000000010000100011",  "000000010000110101",  "000000010001000111",  "000000010001011001",  "000000010001101011",  "000000010001111100",  "000000010010001110",  "000000010010100000",  "000000010010110010",  "000000010011000011",  "000000010011010101",  "000000010011100111",  "000000010011111000",  "000000010100001010",  "000000010100011100",  "000000010100101101",  "000000010100111111",  "000000010101010000",  "000000010101100010",  "000000010101110011",  "000000010110000101",  "000000010110010110",  "000000010110101000",  "000000010110111001",  "000000010111001010",  "000000010111011100",  "000000010111101101",  "000000010111111111",  "000000011000010000",  "000000011000100001",  "000000011000110010",  "000000011001000100",  "000000011001010101",  "000000011001100110",  "000000011001110111",  "000000011010001000",  "000000011010011010",  "000000011010101011",  "000000011010111100",  "000000011011001101",  "000000011011011110",  "000000011011101111",  "000000011100000000",  "000000011100010001",  "000000011100100010",  "000000011100110011",  "000000011101000100",  "000000011101010100",  "000000011101100101",  "000000011101110110",  "000000011110000111",  "000000011110011000",  "000000011110101000",  "000000011110111001",  "000000011111001010",  "000000011111011011",  "000000011111101011",  "000000011111111100",  "000000100000001100",  "000000100000011101",  "000000100000101110",  "000000100000111110",  "000000100001001111",  "000000100001011111",  "000000100001101111",  "000000100010000000",  "000000100010010000",  "000000100010100001",  "000000100010110001",  "000000100011000001",  "000000100011010001",  "000000100011100010",  "000000100011110010",  "000000100100000010",  "000000100100010010",  "000000100100100010",  "000000100100110011",  "000000100101000011",  "000000100101010011",  "000000100101100011",  "000000100101110011",  "000000100110000011",  "000000100110010011",  "000000100110100010",  "000000100110110010",  "000000100111000010",  "000000100111010010",  "000000100111100010",  "000000100111110001",  "000000101000000001",  "000000101000010001",  "000000101000100000",  "000000101000110000",  "000000101001000000",  "000000101001001111",  "000000101001011111",  "000000101001101110",  "000000101001111110",  "000000101010001101",  "000000101010011101",  "000000101010101100",  "000000101010111011",  "000000101011001011",  "000000101011011010",  "000000101011101001",  "000000101011111000",  "000000101100000111",  "000000101100010111",  "000000101100100110",  "000000101100110101",  "000000101101000100",  "000000101101010011",  "000000101101100010",  "000000101101110001",  "000000101110000000",  "000000101110001111",  "000000101110011101",  "000000101110101100",  "000000101110111011",  "000000101111001010",  "000000101111011000",  "000000101111100111",  "000000101111110110",  "000000110000000100",  "000000110000010011",  "000000110000100001",  "000000110000110000",  "000000110000111110",  "000000110001001101",  "000000110001011011",  "000000110001101010",  "000000110001111000",  "000000110010000110",  "000000110010010100",  "000000110010100011",  "000000110010110001",  "000000110010111111",  "000000110011001101",  "000000110011011011",  "000000110011101001",  "000000110011110111",  "000000110100000101",  "000000110100010011",  "000000110100100001",  "000000110100101111",  "000000110100111100",  "000000110101001010",  "000000110101011000",  "000000110101100110",  "000000110101110011",  "000000110110000001",  "000000110110001110",  "000000110110011100",  "000000110110101001",  "000000110110110111",  "000000110111000100",  "000000110111010010",  "000000110111011111",  "000000110111101100",  "000000110111111010",  "000000111000000111",  "000000111000010100",  "000000111000100001",  "000000111000101110",  "000000111000111011",  "000000111001001000",  "000000111001010101",  "000000111001100010",  "000000111001101111",  "000000111001111100",  "000000111010001001",  "000000111010010110",  "000000111010100010",  "000000111010101111",  "000000111010111100",  "000000111011001000",  "000000111011010101",  "000000111011100010",  "000000111011101110",  "000000111011111011",  "000000111100000111",  "000000111100010011",  "000000111100100000",  "000000111100101100",  "000000111100111000",  "000000111101000100",  "000000111101010001",  "000000111101011101",  "000000111101101001",  "000000111101110101",  "000000111110000001",  "000000111110001101",  "000000111110011001",  "000000111110100101",  "000000111110110000",  "000000111110111100",  "000000111111001000",  "000000111111010100",  "000000111111011111",  "000000111111101011",  "000000111111110111",  "000001000000000010",  "000001000000001110",  "000001000000011001",  "000001000000100100",  "000001000000110000",  "000001000000111011",  "000001000001000110",  "000001000001010010",  "000001000001011101",  "000001000001101000",  "000001000001110011",  "000001000001111110",  "000001000010001001",  "000001000010010100",  "000001000010011111",  "000001000010101010",  "000001000010110101",  "000001000010111111",  "000001000011001010",  "000001000011010101",  "000001000011011111",  "000001000011101010",  "000001000011110101",  "000001000011111111",  "000001000100001010",  "000001000100010100",  "000001000100011110",  "000001000100101001",  "000001000100110011",  "000001000100111101",  "000001000101000111",  "000001000101010010",  "000001000101011100",  "000001000101100110",  "000001000101110000",  "000001000101111010",  "000001000110000100",  "000001000110001110",  "000001000110010111",  "000001000110100001",  "000001000110101011",  "000001000110110101",  "000001000110111110",  "000001000111001000",  "000001000111010001",  "000001000111011011",  "000001000111100100",  "000001000111101110",  "000001000111110111",  "000001001000000000",  "000001001000001010",  "000001001000010011",  "000001001000011100",  "000001001000100101",  "000001001000101110",  "000001001000110111",  "000001001001000000",  "000001001001001001",  "000001001001010010",  "000001001001011011",  "000001001001100100",  "000001001001101100",  "000001001001110101",  "000001001001111110",  "000001001010000110",  "000001001010001111",  "000001001010010111",  "000001001010100000",  "000001001010101000",  "000001001010110000",  "000001001010111001",  "000001001011000001",  "000001001011001001",  "000001001011010001",  "000001001011011001",  "000001001011100010",  "000001001011101010",  "000001001011110010",  "000001001011111001",  "000001001100000001",  "000001001100001001",  "000001001100010001",  "000001001100011001",  "000001001100100000",  "000001001100101000",  "000001001100101111",  "000001001100110111",  "000001001100111110",  "000001001101000110",  "000001001101001101",  "000001001101010101",  "000001001101011100",  "000001001101100011",  "000001001101101010",  "000001001101110001",  "000001001101111000",  "000001001101111111",  "000001001110000110",  "000001001110001101",  "000001001110010100",  "000001001110011011",  "000001001110100010",  "000001001110101000",  "000001001110101111",  "000001001110110110",  "000001001110111100",  "000001001111000011",  "000001001111001001",  "000001001111010000",  "000001001111010110",  "000001001111011100",  "000001001111100011",  "000001001111101001",  "000001001111101111",  "000001001111110101",  "000001001111111011",  "000001010000000001",  "000001010000000111",  "000001010000001101",  "000001010000010011",  "000001010000011001",  "000001010000011111",  "000001010000100100",  "000001010000101010",  "000001010000110000",  "000001010000110101",  "000001010000111011",  "000001010001000000",  "000001010001000101",  "000001010001001011",  "000001010001010000",  "000001010001010101",  "000001010001011011",  "000001010001100000",  "000001010001100101",  "000001010001101010",  "000001010001101111",  "000001010001110100",  "000001010001111001",  "000001010001111110",  "000001010010000010",  "000001010010000111",  "000001010010001100",  "000001010010010000",  "000001010010010101",  "000001010010011001",  "000001010010011110",  "000001010010100010",  "000001010010100111",  "000001010010101011",  "000001010010101111",  "000001010010110100",  "000001010010111000",  "000001010010111100",  "000001010011000000",  "000001010011000100",  "000001010011001000",  "000001010011001100",  "000001010011010000",  "000001010011010011",  "000001010011010111",  "000001010011011011",  "000001010011011111",  "000001010011100010",  "000001010011100110",  "000001010011101001",  "000001010011101101",  "000001010011110000",  "000001010011110011",  "000001010011110111",  "000001010011111010",  "000001010011111101",  "000001010100000000",  "000001010100000011",  "000001010100000110",  "000001010100001001",  "000001010100001100",  "000001010100001111",  "000001010100010010",  "000001010100010101",  "000001010100010111",  "000001010100011010",  "000001010100011101",  "000001010100011111",  "000001010100100010",  "000001010100100100",  "000001010100100111",  "000001010100101001",  "000001010100101011",  "000001010100101110",  "000001010100110000",  "000001010100110010",  "000001010100110100",  "000001010100110110",  "000001010100111000",  "000001010100111010",  "000001010100111100",  "000001010100111110",  "000001010100111111",  "000001010101000001",  "000001010101000011",  "000001010101000100",  "000001010101000110",  "000001010101001000",  "000001010101001001",  "000001010101001010",  "000001010101001100",  "000001010101001101",  "000001010101001110",  "000001010101010000",  "000001010101010001",  "000001010101010010",  "000001010101010011",  "000001010101010100",  "000001010101010101",  "000001010101010110",  "000001010101010111",  "000001010101010111",  "000001010101011000",  "000001010101011001",  "000001010101011001",  "000001010101011010",  "000001010101011010",  "000001010101011011",  "000001010101011011",  "000001010101011100",  "000001010101011100",  "000001010101011100",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011101",  "000001010101011100",  "000001010101011100",  "000001010101011100",  "000001010101011100",  "000001010101011011",  "000001010101011011",  "000001010101011010",  "000001010101011010",  "000001010101011001",  "000001010101011000",  "000001010101011000",  "000001010101010111",  "000001010101010110",  "000001010101010101",  "000001010101010100",  "000001010101010011",  "000001010101010010",  "000001010101010001",  "000001010101010000",  "000001010101001111",  "000001010101001110",  "000001010101001101",  "000001010101001011",  "000001010101001010",  "000001010101001000",  "000001010101000111",  "000001010101000101",  "000001010101000100",  "000001010101000010",  "000001010101000001",  "000001010100111111",  "000001010100111101",  "000001010100111011",  "000001010100111001",  "000001010100110111",  "000001010100110110",  "000001010100110011",  "000001010100110001",  "000001010100101111",  "000001010100101101",  "000001010100101011",  "000001010100101001",  "000001010100100110",  "000001010100100100",  "000001010100100001",  "000001010100011111",  "000001010100011100",  "000001010100011010",  "000001010100010111",  "000001010100010101",  "000001010100010010",  "000001010100001111",  "000001010100001100",  "000001010100001001",  "000001010100000110",  "000001010100000011",  "000001010100000000",  "000001010011111101",  "000001010011111010",  "000001010011110111",  "000001010011110100",  "000001010011110000",  "000001010011101101",  "000001010011101010",  "000001010011100110",  "000001010011100011",  "000001010011011111",  "000001010011011100",  "000001010011011000",  "000001010011010101",  "000001010011010001",  "000001010011001101",  "000001010011001001",  "000001010011000101",  "000001010011000001",  "000001010010111101",  "000001010010111001",  "000001010010110101",  "000001010010110001",  "000001010010101101",  "000001010010101001",  "000001010010100101",  "000001010010100000",  "000001010010011100",  "000001010010011000",  "000001010010010011",  "000001010010001111",  "000001010010001010",  "000001010010000110",  "000001010010000001",  "000001010001111100",  "000001010001111000",  "000001010001110011",  "000001010001101110",  "000001010001101001",  "000001010001100100",  "000001010001011111",  "000001010001011010",  "000001010001010101",  "000001010001010000",  "000001010001001011",  "000001010001000110",  "000001010001000000",  "000001010000111011",  "000001010000110110",  "000001010000110000",  "000001010000101011",  "000001010000100101",  "000001010000100000",  "000001010000011010",  "000001010000010101",  "000001010000001111",  "000001010000001001",  "000001010000000100",  "000001001111111110",  "000001001111111000",  "000001001111110010",  "000001001111101100",  "000001001111100110",  "000001001111100000",  "000001001111011010",  "000001001111010100",  "000001001111001110",  "000001001111000111",  "000001001111000001",  "000001001110111011",  "000001001110110100",  "000001001110101110",  "000001001110101000",  "000001001110100001",  "000001001110011011",  "000001001110010100",  "000001001110001101",  "000001001110000111",  "000001001110000000",  "000001001101111001",  "000001001101110010",  "000001001101101100",  "000001001101100101",  "000001001101011110",  "000001001101010111",  "000001001101010000",  "000001001101001001",  "000001001101000010",  "000001001100111010",  "000001001100110011",  "000001001100101100",  "000001001100100101",  "000001001100011101",  "000001001100010110",  "000001001100001111",  "000001001100000111",  "000001001100000000",  "000001001011111000",  "000001001011110001",  "000001001011101001",  "000001001011100001",  "000001001011011010",  "000001001011010010",  "000001001011001010",  "000001001011000010",  "000001001010111010",  "000001001010110010",  "000001001010101010",  "000001001010100010",  "000001001010011010",  "000001001010010010",  "000001001010001010",  "000001001010000010",  "000001001001111010",  "000001001001110001",  "000001001001101001",  "000001001001100001",  "000001001001011000",  "000001001001010000",  "000001001001001000",  "000001001000111111",  "000001001000110110",  "000001001000101110",  "000001001000100101",  "000001001000011101",  "000001001000010100",  "000001001000001011",  "000001001000000010",  "000001000111111010",  "000001000111110001",  "000001000111101000",  "000001000111011111",  "000001000111010110",  "000001000111001101",  "000001000111000100",  "000001000110111011",  "000001000110110001",  "000001000110101000",  "000001000110011111",  "000001000110010110",  "000001000110001101",  "000001000110000011",  "000001000101111010",  "000001000101110000",  "000001000101100111",  "000001000101011101",  "000001000101010100",  "000001000101001010",  "000001000101000001",  "000001000100110111",  "000001000100101101",  "000001000100100100",  "000001000100011010",  "000001000100010000",  "000001000100000110",  "000001000011111100",  "000001000011110010",  "000001000011101001",  "000001000011011111",  "000001000011010101",  "000001000011001010",  "000001000011000000",  "000001000010110110",  "000001000010101100",  "000001000010100010",  "000001000010011000",  "000001000010001101",  "000001000010000011",  "000001000001111001",  "000001000001101110",  "000001000001100100",  "000001000001011001",  "000001000001001111",  "000001000001000100",  "000001000000111010",  "000001000000101111",  "000001000000100101",  "000001000000011010",  "000001000000001111",  "000001000000000101",  "000000111111111010",  "000000111111101111",  "000000111111100100",  "000000111111011001",  "000000111111001110",  "000000111111000100",  "000000111110111001",  "000000111110101110",  "000000111110100010",  "000000111110010111",  "000000111110001100",  "000000111110000001",  "000000111101110110",  "000000111101101011",  "000000111101100000",  "000000111101010100",  "000000111101001001",  "000000111100111110",  "000000111100110010",  "000000111100100111",  "000000111100011011",  "000000111100010000",  "000000111100000101",  "000000111011111001",  "000000111011101101",  "000000111011100010",  "000000111011010110",  "000000111011001011",  "000000111010111111",  "000000111010110011",  "000000111010100111",  "000000111010011100",  "000000111010010000",  "000000111010000100",  "000000111001111000",  "000000111001101100",  "000000111001100000",  "000000111001010100",  "000000111001001000",  "000000111000111100",  "000000111000110000",  "000000111000100100",  "000000111000011000",  "000000111000001100",  "000000111000000000",  "000000110111110100",  "000000110111100111",  "000000110111011011",  "000000110111001111",  "000000110111000011",  "000000110110110110",  "000000110110101010",  "000000110110011101",  "000000110110010001",  "000000110110000101",  "000000110101111000",  "000000110101101100",  "000000110101011111",  "000000110101010010",  "000000110101000110",  "000000110100111001",  "000000110100101101",  "000000110100100000",  "000000110100010011",  "000000110100000111",  "000000110011111010",  "000000110011101101",  "000000110011100000",  "000000110011010011",  "000000110011000111",  "000000110010111010",  "000000110010101101",  "000000110010100000",  "000000110010010011",  "000000110010000110",  "000000110001111001",  "000000110001101100",  "000000110001011111",  "000000110001010010",  "000000110001000101",  "000000110000110111",  "000000110000101010",  "000000110000011101",  "000000110000010000",  "000000110000000011",  "000000101111110101",  "000000101111101000",  "000000101111011011",  "000000101111001110",  "000000101111000000",  "000000101110110011",  "000000101110100101",  "000000101110011000",  "000000101110001011",  "000000101101111101",  "000000101101110000",  "000000101101100010",  "000000101101010101",  "000000101101000111",  "000000101100111010",  "000000101100101100",  "000000101100011110",  "000000101100010001",  "000000101100000011",  "000000101011110101",  "000000101011101000",  "000000101011011010",  "000000101011001100",  "000000101010111110",  "000000101010110001",  "000000101010100011",  "000000101010010101",  "000000101010000111",  "000000101001111001",  "000000101001101011",  "000000101001011110",  "000000101001010000",  "000000101001000010",  "000000101000110100",  "000000101000100110",  "000000101000011000",  "000000101000001010",  "000000100111111100",  "000000100111101110",  "000000100111100000",  "000000100111010001",  "000000100111000011",  "000000100110110101",  "000000100110100111",  "000000100110011001",  "000000100110001011",  "000000100101111100",  "000000100101101110",  "000000100101100000",  "000000100101010010",  "000000100101000100",  "000000100100110101",  "000000100100100111",  "000000100100011001",  "000000100100001010",  "000000100011111100",  "000000100011101110",  "000000100011011111",  "000000100011010001",  "000000100011000010",  "000000100010110100",  "000000100010100101",  "000000100010010111",  "000000100010001001",  "000000100001111010",  "000000100001101100",  "000000100001011101",  "000000100001001110",  "000000100001000000",  "000000100000110001",  "000000100000100011",  "000000100000010100",  "000000100000000110",  "000000011111110111",  "000000011111101000",  "000000011111011010",  "000000011111001011",  "000000011110111100",  "000000011110101110",  "000000011110011111",  "000000011110010000",  "000000011110000010",  "000000011101110011",  "000000011101100100",  "000000011101010101",  "000000011101000111",  "000000011100111000",  "000000011100101001",  "000000011100011010",  "000000011100001011",  "000000011011111100",  "000000011011101110",  "000000011011011111",  "000000011011010000",  "000000011011000001",  "000000011010110010",  "000000011010100011",  "000000011010010100",  "000000011010000101",  "000000011001110111",  "000000011001101000",  "000000011001011001",  "000000011001001010",  "000000011000111011",  "000000011000101100",  "000000011000011101",  "000000011000001110",  "000000010111111111",  "000000010111110000",  "000000010111100001",  "000000010111010010",  "000000010111000011",  "000000010110110100",  "000000010110100101",  "000000010110010110",  "000000010110000110",  "000000010101110111",  "000000010101101000",  "000000010101011001",  "000000010101001010",  "000000010100111011",  "000000010100101100",  "000000010100011101",  "000000010100001110",  "000000010011111111",  "000000010011101111",  "000000010011100000",  "000000010011010001",  "000000010011000010",  "000000010010110011",  "000000010010100100",  "000000010010010101",  "000000010010000101",  "000000010001110110",  "000000010001100111",  "000000010001011000",  "000000010001001001",  "000000010000111001",  "000000010000101010",  "000000010000011011",  "000000010000001100",  "000000001111111101",  "000000001111101101",  "000000001111011110",  "000000001111001111",  "000000001111000000",  "000000001110110000",  "000000001110100001",  "000000001110010010",  "000000001110000011",  "000000001101110100",  "000000001101100100",  "000000001101010101",  "000000001101000110",  "000000001100110111",  "000000001100100111",  "000000001100011000",  "000000001100001001",  "000000001011111001",  "000000001011101010",  "000000001011011011",  "000000001011001100",  "000000001010111100",  "000000001010101101",  "000000001010011110",  "000000001010001111",  "000000001001111111",  "000000001001110000",  "000000001001100001",  "000000001001010010",  "000000001001000010",  "000000001000110011",  "000000001000100100",  "000000001000010101",  "000000001000000101",  "000000000111110110",  "000000000111100111",  "000000000111011000",  "000000000111001000",  "000000000110111001",  "000000000110101010",  "000000000110011011",  "000000000110001011",  "000000000101111100",  "000000000101101101",  "000000000101011110",  "000000000101001110",  "000000000100111111",  "000000000100110000",  "000000000100100001",  "000000000100010001",  "000000000100000010",  "000000000011110011",  "000000000011100100",  "000000000011010101",  "000000000011000101",  "000000000010110110",  "000000000010100111",  "000000000010011000",  "000000000010001001",  "000000000001111001",  "000000000001101010",  "000000000001011011",  "000000000001001100",  "000000000000111101",  "000000000000101101",  "000000000000011110",  "000000000000001111"),("000000000000000000",  "111111111111110001",  "111111111111100010",  "111111111111010011",  "111111111111000011",  "111111111110110100",  "111111111110100101",  "111111111110010110",  "111111111110000111",  "111111111101111000",  "111111111101101001",  "111111111101011010",  "111111111101001011",  "111111111100111100",  "111111111100101101",  "111111111100011110",  "111111111100001111",  "111111111100000000",  "111111111011110001",  "111111111011100010",  "111111111011010010",  "111111111011000100",  "111111111010110101",  "111111111010100110",  "111111111010010111",  "111111111010001000",  "111111111001111001",  "111111111001101010",  "111111111001011011",  "111111111001001100",  "111111111000111101",  "111111111000101110",  "111111111000011111",  "111111111000010000",  "111111111000000001",  "111111110111110011",  "111111110111100100",  "111111110111010101",  "111111110111000110",  "111111110110110111",  "111111110110101000",  "111111110110011010",  "111111110110001011",  "111111110101111100",  "111111110101101101",  "111111110101011111",  "111111110101010000",  "111111110101000001",  "111111110100110010",  "111111110100100100",  "111111110100010101",  "111111110100000110",  "111111110011111000",  "111111110011101001",  "111111110011011010",  "111111110011001100",  "111111110010111101",  "111111110010101111",  "111111110010100000",  "111111110010010001",  "111111110010000011",  "111111110001110100",  "111111110001100110",  "111111110001010111",  "111111110001001001",  "111111110000111010",  "111111110000101100",  "111111110000011101",  "111111110000001111",  "111111110000000001",  "111111101111110010",  "111111101111100100",  "111111101111010101",  "111111101111000111",  "111111101110111001",  "111111101110101010",  "111111101110011100",  "111111101110001110",  "111111101110000000",  "111111101101110001",  "111111101101100011",  "111111101101010101",  "111111101101000111",  "111111101100111000",  "111111101100101010",  "111111101100011100",  "111111101100001110",  "111111101100000000",  "111111101011110010",  "111111101011100100",  "111111101011010110",  "111111101011000111",  "111111101010111001",  "111111101010101011",  "111111101010011101",  "111111101010001111",  "111111101010000001",  "111111101001110011",  "111111101001100110",  "111111101001011000",  "111111101001001010",  "111111101000111100",  "111111101000101110",  "111111101000100000",  "111111101000010010",  "111111101000000101",  "111111100111110111",  "111111100111101001",  "111111100111011011",  "111111100111001110",  "111111100111000000",  "111111100110110010",  "111111100110100101",  "111111100110010111",  "111111100110001001",  "111111100101111100",  "111111100101101110",  "111111100101100001",  "111111100101010011",  "111111100101000110",  "111111100100111000",  "111111100100101011",  "111111100100011101",  "111111100100010000",  "111111100100000010",  "111111100011110101",  "111111100011101000",  "111111100011011010",  "111111100011001101",  "111111100011000000",  "111111100010110011",  "111111100010100101",  "111111100010011000",  "111111100010001011",  "111111100001111110",  "111111100001110001",  "111111100001100011",  "111111100001010110",  "111111100001001001",  "111111100000111100",  "111111100000101111",  "111111100000100010",  "111111100000010101",  "111111100000001000",  "111111011111111011",  "111111011111101110",  "111111011111100001",  "111111011111010101",  "111111011111001000",  "111111011110111011",  "111111011110101110",  "111111011110100001",  "111111011110010101",  "111111011110001000",  "111111011101111011",  "111111011101101111",  "111111011101100010",  "111111011101010101",  "111111011101001001",  "111111011100111100",  "111111011100110000",  "111111011100100011",  "111111011100010111",  "111111011100001010",  "111111011011111110",  "111111011011110001",  "111111011011100101",  "111111011011011001",  "111111011011001100",  "111111011011000000",  "111111011010110100",  "111111011010101000",  "111111011010011011",  "111111011010001111",  "111111011010000011",  "111111011001110111",  "111111011001101011",  "111111011001011111",  "111111011001010011",  "111111011001000111",  "111111011000111011",  "111111011000101111",  "111111011000100011",  "111111011000010111",  "111111011000001011",  "111111010111111111",  "111111010111110011",  "111111010111101000",  "111111010111011100",  "111111010111010000",  "111111010111000100",  "111111010110111001",  "111111010110101101",  "111111010110100001",  "111111010110010110",  "111111010110001010",  "111111010101111111",  "111111010101110011",  "111111010101101000",  "111111010101011100",  "111111010101010001",  "111111010101000110",  "111111010100111010",  "111111010100101111",  "111111010100100100",  "111111010100011000",  "111111010100001101",  "111111010100000010",  "111111010011110111",  "111111010011101100",  "111111010011100001",  "111111010011010101",  "111111010011001010",  "111111010010111111",  "111111010010110100",  "111111010010101001",  "111111010010011111",  "111111010010010100",  "111111010010001001",  "111111010001111110",  "111111010001110011",  "111111010001101000",  "111111010001011110",  "111111010001010011",  "111111010001001000",  "111111010000111110",  "111111010000110011",  "111111010000101001",  "111111010000011110",  "111111010000010100",  "111111010000001001",  "111111001111111111",  "111111001111110100",  "111111001111101010",  "111111001111100000",  "111111001111010101",  "111111001111001011",  "111111001111000001",  "111111001110110111",  "111111001110101100",  "111111001110100010",  "111111001110011000",  "111111001110001110",  "111111001110000100",  "111111001101111010",  "111111001101110000",  "111111001101100110",  "111111001101011100",  "111111001101010011",  "111111001101001001",  "111111001100111111",  "111111001100110101",  "111111001100101011",  "111111001100100010",  "111111001100011000",  "111111001100001110",  "111111001100000101",  "111111001011111011",  "111111001011110010",  "111111001011101000",  "111111001011011111",  "111111001011010110",  "111111001011001100",  "111111001011000011",  "111111001010111010",  "111111001010110000",  "111111001010100111",  "111111001010011110",  "111111001010010101",  "111111001010001100",  "111111001010000010",  "111111001001111001",  "111111001001110000",  "111111001001100111",  "111111001001011110",  "111111001001010110",  "111111001001001101",  "111111001001000100",  "111111001000111011",  "111111001000110010",  "111111001000101010",  "111111001000100001",  "111111001000011000",  "111111001000010000",  "111111001000000111",  "111111000111111111",  "111111000111110110",  "111111000111101110",  "111111000111100101",  "111111000111011101",  "111111000111010100",  "111111000111001100",  "111111000111000100",  "111111000110111100",  "111111000110110011",  "111111000110101011",  "111111000110100011",  "111111000110011011",  "111111000110010011",  "111111000110001011",  "111111000110000011",  "111111000101111011",  "111111000101110011",  "111111000101101011",  "111111000101100100",  "111111000101011100",  "111111000101010100",  "111111000101001100",  "111111000101000101",  "111111000100111101",  "111111000100110101",  "111111000100101110",  "111111000100100110",  "111111000100011111",  "111111000100010111",  "111111000100010000",  "111111000100001001",  "111111000100000001",  "111111000011111010",  "111111000011110011",  "111111000011101100",  "111111000011100100",  "111111000011011101",  "111111000011010110",  "111111000011001111",  "111111000011001000",  "111111000011000001",  "111111000010111010",  "111111000010110011",  "111111000010101101",  "111111000010100110",  "111111000010011111",  "111111000010011000",  "111111000010010010",  "111111000010001011",  "111111000010000100",  "111111000001111110",  "111111000001110111",  "111111000001110001",  "111111000001101010",  "111111000001100100",  "111111000001011110",  "111111000001010111",  "111111000001010001",  "111111000001001011",  "111111000001000100",  "111111000000111110",  "111111000000111000",  "111111000000110010",  "111111000000101100",  "111111000000100110",  "111111000000100000",  "111111000000011010",  "111111000000010100",  "111111000000001110",  "111111000000001001",  "111111000000000011",  "111110111111111101",  "111110111111110111",  "111110111111110010",  "111110111111101100",  "111110111111100111",  "111110111111100001",  "111110111111011100",  "111110111111010110",  "111110111111010001",  "111110111111001011",  "111110111111000110",  "111110111111000001",  "111110111110111100",  "111110111110110110",  "111110111110110001",  "111110111110101100",  "111110111110100111",  "111110111110100010",  "111110111110011101",  "111110111110011000",  "111110111110010011",  "111110111110001110",  "111110111110001010",  "111110111110000101",  "111110111110000000",  "111110111101111011",  "111110111101110111",  "111110111101110010",  "111110111101101110",  "111110111101101001",  "111110111101100101",  "111110111101100000",  "111110111101011100",  "111110111101010111",  "111110111101010011",  "111110111101001111",  "111110111101001011",  "111110111101000110",  "111110111101000010",  "111110111100111110",  "111110111100111010",  "111110111100110110",  "111110111100110010",  "111110111100101110",  "111110111100101010",  "111110111100100110",  "111110111100100011",  "111110111100011111",  "111110111100011011",  "111110111100010111",  "111110111100010100",  "111110111100010000",  "111110111100001101",  "111110111100001001",  "111110111100000110",  "111110111100000010",  "111110111011111111",  "111110111011111100",  "111110111011111000",  "111110111011110101",  "111110111011110010",  "111110111011101111",  "111110111011101011",  "111110111011101000",  "111110111011100101",  "111110111011100010",  "111110111011011111",  "111110111011011100",  "111110111011011010",  "111110111011010111",  "111110111011010100",  "111110111011010001",  "111110111011001111",  "111110111011001100",  "111110111011001001",  "111110111011000111",  "111110111011000100",  "111110111011000010",  "111110111010111111",  "111110111010111101",  "111110111010111010",  "111110111010111000",  "111110111010110110",  "111110111010110100",  "111110111010110001",  "111110111010101111",  "111110111010101101",  "111110111010101011",  "111110111010101001",  "111110111010100111",  "111110111010100101",  "111110111010100011",  "111110111010100001",  "111110111010100000",  "111110111010011110",  "111110111010011100",  "111110111010011010",  "111110111010011001",  "111110111010010111",  "111110111010010110",  "111110111010010100",  "111110111010010011",  "111110111010010001",  "111110111010010000",  "111110111010001110",  "111110111010001101",  "111110111010001100",  "111110111010001011",  "111110111010001001",  "111110111010001000",  "111110111010000111",  "111110111010000110",  "111110111010000101",  "111110111010000100",  "111110111010000011",  "111110111010000010",  "111110111010000010",  "111110111010000001",  "111110111010000000",  "111110111001111111",  "111110111001111111",  "111110111001111110",  "111110111001111110",  "111110111001111101",  "111110111001111101",  "111110111001111100",  "111110111001111100",  "111110111001111011",  "111110111001111011",  "111110111001111011",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111010",  "111110111001111011",  "111110111001111011",  "111110111001111011",  "111110111001111100",  "111110111001111100",  "111110111001111100",  "111110111001111101",  "111110111001111101",  "111110111001111110",  "111110111001111111",  "111110111001111111",  "111110111010000000",  "111110111010000001",  "111110111010000001",  "111110111010000010",  "111110111010000011",  "111110111010000100",  "111110111010000101",  "111110111010000110",  "111110111010000111",  "111110111010001000",  "111110111010001001",  "111110111010001010",  "111110111010001100",  "111110111010001101",  "111110111010001110",  "111110111010001111",  "111110111010010001",  "111110111010010010",  "111110111010010100",  "111110111010010101",  "111110111010010111",  "111110111010011000",  "111110111010011010",  "111110111010011011",  "111110111010011101",  "111110111010011111",  "111110111010100001",  "111110111010100011",  "111110111010100100",  "111110111010100110",  "111110111010101000",  "111110111010101010",  "111110111010101100",  "111110111010101110",  "111110111010110000",  "111110111010110011",  "111110111010110101",  "111110111010110111",  "111110111010111001",  "111110111010111100",  "111110111010111110",  "111110111011000000",  "111110111011000011",  "111110111011000101",  "111110111011001000",  "111110111011001010",  "111110111011001101",  "111110111011010000",  "111110111011010010",  "111110111011010101",  "111110111011011000",  "111110111011011010",  "111110111011011101",  "111110111011100000",  "111110111011100011",  "111110111011100110",  "111110111011101001",  "111110111011101100",  "111110111011101111",  "111110111011110010",  "111110111011110101",  "111110111011111001",  "111110111011111100",  "111110111011111111",  "111110111100000011",  "111110111100000110",  "111110111100001001",  "111110111100001101",  "111110111100010000",  "111110111100010100",  "111110111100010111",  "111110111100011011",  "111110111100011111",  "111110111100100010",  "111110111100100110",  "111110111100101010",  "111110111100101101",  "111110111100110001",  "111110111100110101",  "111110111100111001",  "111110111100111101",  "111110111101000001",  "111110111101000101",  "111110111101001001",  "111110111101001101",  "111110111101010001",  "111110111101010110",  "111110111101011010",  "111110111101011110",  "111110111101100010",  "111110111101100111",  "111110111101101011",  "111110111101101111",  "111110111101110100",  "111110111101111000",  "111110111101111101",  "111110111110000010",  "111110111110000110",  "111110111110001011",  "111110111110001111",  "111110111110010100",  "111110111110011001",  "111110111110011110",  "111110111110100011",  "111110111110100111",  "111110111110101100",  "111110111110110001",  "111110111110110110",  "111110111110111011",  "111110111111000000",  "111110111111000101",  "111110111111001011",  "111110111111010000",  "111110111111010101",  "111110111111011010",  "111110111111100000",  "111110111111100101",  "111110111111101010",  "111110111111110000",  "111110111111110101",  "111110111111111011",  "111111000000000000",  "111111000000000110",  "111111000000001011",  "111111000000010001",  "111111000000010110",  "111111000000011100",  "111111000000100010",  "111111000000101000",  "111111000000101101",  "111111000000110011",  "111111000000111001",  "111111000000111111",  "111111000001000101",  "111111000001001011",  "111111000001010001",  "111111000001010111",  "111111000001011101",  "111111000001100011",  "111111000001101001",  "111111000001110000",  "111111000001110110",  "111111000001111100",  "111111000010000010",  "111111000010001001",  "111111000010001111",  "111111000010010101",  "111111000010011100",  "111111000010100010",  "111111000010101001",  "111111000010101111",  "111111000010110110",  "111111000010111101",  "111111000011000011",  "111111000011001010",  "111111000011010001",  "111111000011010111",  "111111000011011110",  "111111000011100101",  "111111000011101100",  "111111000011110011",  "111111000011111010",  "111111000100000000",  "111111000100000111",  "111111000100001110",  "111111000100010110",  "111111000100011101",  "111111000100100100",  "111111000100101011",  "111111000100110010",  "111111000100111001",  "111111000101000001",  "111111000101001000",  "111111000101001111",  "111111000101010110",  "111111000101011110",  "111111000101100101",  "111111000101101101",  "111111000101110100",  "111111000101111100",  "111111000110000011",  "111111000110001011",  "111111000110010010",  "111111000110011010",  "111111000110100010",  "111111000110101001",  "111111000110110001",  "111111000110111001",  "111111000111000001",  "111111000111001001",  "111111000111010000",  "111111000111011000",  "111111000111100000",  "111111000111101000",  "111111000111110000",  "111111000111111000",  "111111001000000000",  "111111001000001000",  "111111001000010000",  "111111001000011001",  "111111001000100001",  "111111001000101001",  "111111001000110001",  "111111001000111001",  "111111001001000010",  "111111001001001010",  "111111001001010010",  "111111001001011011",  "111111001001100011",  "111111001001101100",  "111111001001110100",  "111111001001111101",  "111111001010000101",  "111111001010001110",  "111111001010010110",  "111111001010011111",  "111111001010101000",  "111111001010110000",  "111111001010111001",  "111111001011000010",  "111111001011001010",  "111111001011010011",  "111111001011011100",  "111111001011100101",  "111111001011101110",  "111111001011110111",  "111111001100000000",  "111111001100001001",  "111111001100010010",  "111111001100011011",  "111111001100100100",  "111111001100101101",  "111111001100110110",  "111111001100111111",  "111111001101001000",  "111111001101010001",  "111111001101011010",  "111111001101100100",  "111111001101101101",  "111111001101110110",  "111111001110000000",  "111111001110001001",  "111111001110010010",  "111111001110011100",  "111111001110100101",  "111111001110101111",  "111111001110111000",  "111111001111000001",  "111111001111001011",  "111111001111010101",  "111111001111011110",  "111111001111101000",  "111111001111110001",  "111111001111111011",  "111111010000000101",  "111111010000001110",  "111111010000011000",  "111111010000100010",  "111111010000101100",  "111111010000110110",  "111111010000111111",  "111111010001001001",  "111111010001010011",  "111111010001011101",  "111111010001100111",  "111111010001110001",  "111111010001111011",  "111111010010000101",  "111111010010001111",  "111111010010011001",  "111111010010100011",  "111111010010101101",  "111111010010110111",  "111111010011000001",  "111111010011001100",  "111111010011010110",  "111111010011100000",  "111111010011101010",  "111111010011110100",  "111111010011111111",  "111111010100001001",  "111111010100010011",  "111111010100011110",  "111111010100101000",  "111111010100110011",  "111111010100111101",  "111111010101000111",  "111111010101010010",  "111111010101011100",  "111111010101100111",  "111111010101110001",  "111111010101111100",  "111111010110000111",  "111111010110010001",  "111111010110011100",  "111111010110100110",  "111111010110110001",  "111111010110111100",  "111111010111000110",  "111111010111010001",  "111111010111011100",  "111111010111100111",  "111111010111110001",  "111111010111111100",  "111111011000000111",  "111111011000010010",  "111111011000011101",  "111111011000101000",  "111111011000110011",  "111111011000111101",  "111111011001001000",  "111111011001010011",  "111111011001011110",  "111111011001101001",  "111111011001110100",  "111111011001111111",  "111111011010001010",  "111111011010010110",  "111111011010100001",  "111111011010101100",  "111111011010110111",  "111111011011000010",  "111111011011001101",  "111111011011011000",  "111111011011100100",  "111111011011101111",  "111111011011111010",  "111111011100000101",  "111111011100010001",  "111111011100011100",  "111111011100100111",  "111111011100110010",  "111111011100111110",  "111111011101001001",  "111111011101010101",  "111111011101100000",  "111111011101101011",  "111111011101110111",  "111111011110000010",  "111111011110001110",  "111111011110011001",  "111111011110100101",  "111111011110110000",  "111111011110111100",  "111111011111000111",  "111111011111010011",  "111111011111011110",  "111111011111101010",  "111111011111110110",  "111111100000000001",  "111111100000001101",  "111111100000011000",  "111111100000100100",  "111111100000110000",  "111111100000111011",  "111111100001000111",  "111111100001010011",  "111111100001011111",  "111111100001101010",  "111111100001110110",  "111111100010000010",  "111111100010001110",  "111111100010011010",  "111111100010100101",  "111111100010110001",  "111111100010111101",  "111111100011001001",  "111111100011010101",  "111111100011100001",  "111111100011101100",  "111111100011111000",  "111111100100000100",  "111111100100010000",  "111111100100011100",  "111111100100101000",  "111111100100110100",  "111111100101000000",  "111111100101001100",  "111111100101011000",  "111111100101100100",  "111111100101110000",  "111111100101111100",  "111111100110001000",  "111111100110010100",  "111111100110100000",  "111111100110101100",  "111111100110111001",  "111111100111000101",  "111111100111010001",  "111111100111011101",  "111111100111101001",  "111111100111110101",  "111111101000000001",  "111111101000001110",  "111111101000011010",  "111111101000100110",  "111111101000110010",  "111111101000111110",  "111111101001001010",  "111111101001010111",  "111111101001100011",  "111111101001101111",  "111111101001111011",  "111111101010001000",  "111111101010010100",  "111111101010100000",  "111111101010101101",  "111111101010111001",  "111111101011000101",  "111111101011010001",  "111111101011011110",  "111111101011101010",  "111111101011110110",  "111111101100000011",  "111111101100001111",  "111111101100011011",  "111111101100101000",  "111111101100110100",  "111111101101000001",  "111111101101001101",  "111111101101011001",  "111111101101100110",  "111111101101110010",  "111111101101111111",  "111111101110001011",  "111111101110010111",  "111111101110100100",  "111111101110110000",  "111111101110111101",  "111111101111001001",  "111111101111010110",  "111111101111100010",  "111111101111101111",  "111111101111111011",  "111111110000001000",  "111111110000010100",  "111111110000100000",  "111111110000101101",  "111111110000111001",  "111111110001000110",  "111111110001010010",  "111111110001011111",  "111111110001101011",  "111111110001111000",  "111111110010000101",  "111111110010010001",  "111111110010011110",  "111111110010101010",  "111111110010110111",  "111111110011000011",  "111111110011010000",  "111111110011011100",  "111111110011101001",  "111111110011110101",  "111111110100000010",  "111111110100001110",  "111111110100011011",  "111111110100101000",  "111111110100110100",  "111111110101000001",  "111111110101001101",  "111111110101011010",  "111111110101100110",  "111111110101110011",  "111111110110000000",  "111111110110001100",  "111111110110011001",  "111111110110100101",  "111111110110110010",  "111111110110111110",  "111111110111001011",  "111111110111011000",  "111111110111100100",  "111111110111110001",  "111111110111111101",  "111111111000001010",  "111111111000010110",  "111111111000100011",  "111111111000110000",  "111111111000111100",  "111111111001001001",  "111111111001010101",  "111111111001100010",  "111111111001101111",  "111111111001111011",  "111111111010001000",  "111111111010010100",  "111111111010100001",  "111111111010101101",  "111111111010111010",  "111111111011000111",  "111111111011010011",  "111111111011100000",  "111111111011101100",  "111111111011111001",  "111111111100000101",  "111111111100010010",  "111111111100011111",  "111111111100101011",  "111111111100111000",  "111111111101000100",  "111111111101010001",  "111111111101011101",  "111111111101101010",  "111111111101110110",  "111111111110000011",  "111111111110001111",  "111111111110011100",  "111111111110101000",  "111111111110110101",  "111111111111000001",  "111111111111001110",  "111111111111011011",  "111111111111100111",  "111111111111110100"),("000000000000000000",  "000000000000001100",  "000000000000011001",  "000000000000100101",  "000000000000110010",  "000000000000111110",  "000000000001001011",  "000000000001010111",  "000000000001100100",  "000000000001110000",  "000000000001111101",  "000000000010001001",  "000000000010010110",  "000000000010100010",  "000000000010101110",  "000000000010111011",  "000000000011000111",  "000000000011010100",  "000000000011100000",  "000000000011101100",  "000000000011111001",  "000000000100000101",  "000000000100010010",  "000000000100011110",  "000000000100101010",  "000000000100110111",  "000000000101000011",  "000000000101001111",  "000000000101011100",  "000000000101101000",  "000000000101110100",  "000000000110000000",  "000000000110001101",  "000000000110011001",  "000000000110100101",  "000000000110110010",  "000000000110111110",  "000000000111001010",  "000000000111010110",  "000000000111100011",  "000000000111101111",  "000000000111111011",  "000000001000000111",  "000000001000010011",  "000000001000100000",  "000000001000101100",  "000000001000111000",  "000000001001000100",  "000000001001010000",  "000000001001011100",  "000000001001101000",  "000000001001110101",  "000000001010000001",  "000000001010001101",  "000000001010011001",  "000000001010100101",  "000000001010110001",  "000000001010111101",  "000000001011001001",  "000000001011010101",  "000000001011100001",  "000000001011101101",  "000000001011111001",  "000000001100000101",  "000000001100010001",  "000000001100011101",  "000000001100101001",  "000000001100110101",  "000000001101000001",  "000000001101001101",  "000000001101011001",  "000000001101100101",  "000000001101110000",  "000000001101111100",  "000000001110001000",  "000000001110010100",  "000000001110100000",  "000000001110101100",  "000000001110110111",  "000000001111000011",  "000000001111001111",  "000000001111011011",  "000000001111100110",  "000000001111110010",  "000000001111111110",  "000000010000001010",  "000000010000010101",  "000000010000100001",  "000000010000101101",  "000000010000111000",  "000000010001000100",  "000000010001001111",  "000000010001011011",  "000000010001100111",  "000000010001110010",  "000000010001111110",  "000000010010001001",  "000000010010010101",  "000000010010100000",  "000000010010101100",  "000000010010110111",  "000000010011000011",  "000000010011001110",  "000000010011011010",  "000000010011100101",  "000000010011110000",  "000000010011111100",  "000000010100000111",  "000000010100010011",  "000000010100011110",  "000000010100101001",  "000000010100110101",  "000000010101000000",  "000000010101001011",  "000000010101010110",  "000000010101100010",  "000000010101101101",  "000000010101111000",  "000000010110000011",  "000000010110001110",  "000000010110011010",  "000000010110100101",  "000000010110110000",  "000000010110111011",  "000000010111000110",  "000000010111010001",  "000000010111011100",  "000000010111100111",  "000000010111110010",  "000000010111111101",  "000000011000001000",  "000000011000010011",  "000000011000011110",  "000000011000101001",  "000000011000110100",  "000000011000111111",  "000000011001001001",  "000000011001010100",  "000000011001011111",  "000000011001101010",  "000000011001110101",  "000000011001111111",  "000000011010001010",  "000000011010010101",  "000000011010100000",  "000000011010101010",  "000000011010110101",  "000000011011000000",  "000000011011001010",  "000000011011010101",  "000000011011011111",  "000000011011101010",  "000000011011110100",  "000000011011111111",  "000000011100001001",  "000000011100010100",  "000000011100011110",  "000000011100101001",  "000000011100110011",  "000000011100111110",  "000000011101001000",  "000000011101010010",  "000000011101011101",  "000000011101100111",  "000000011101110001",  "000000011101111011",  "000000011110000110",  "000000011110010000",  "000000011110011010",  "000000011110100100",  "000000011110101110",  "000000011110111001",  "000000011111000011",  "000000011111001101",  "000000011111010111",  "000000011111100001",  "000000011111101011",  "000000011111110101",  "000000011111111111",  "000000100000001001",  "000000100000010011",  "000000100000011101",  "000000100000100111",  "000000100000110000",  "000000100000111010",  "000000100001000100",  "000000100001001110",  "000000100001011000",  "000000100001100001",  "000000100001101011",  "000000100001110101",  "000000100001111110",  "000000100010001000",  "000000100010010010",  "000000100010011011",  "000000100010100101",  "000000100010101110",  "000000100010111000",  "000000100011000001",  "000000100011001011",  "000000100011010100",  "000000100011011110",  "000000100011100111",  "000000100011110000",  "000000100011111010",  "000000100100000011",  "000000100100001100",  "000000100100010110",  "000000100100011111",  "000000100100101000",  "000000100100110001",  "000000100100111011",  "000000100101000100",  "000000100101001101",  "000000100101010110",  "000000100101011111",  "000000100101101000",  "000000100101110001",  "000000100101111010",  "000000100110000011",  "000000100110001100",  "000000100110010101",  "000000100110011110",  "000000100110100111",  "000000100110101111",  "000000100110111000",  "000000100111000001",  "000000100111001010",  "000000100111010010",  "000000100111011011",  "000000100111100100",  "000000100111101100",  "000000100111110101",  "000000100111111110",  "000000101000000110",  "000000101000001111",  "000000101000010111",  "000000101000100000",  "000000101000101000",  "000000101000110001",  "000000101000111001",  "000000101001000001",  "000000101001001010",  "000000101001010010",  "000000101001011010",  "000000101001100011",  "000000101001101011",  "000000101001110011",  "000000101001111011",  "000000101010000011",  "000000101010001011",  "000000101010010011",  "000000101010011100",  "000000101010100100",  "000000101010101100",  "000000101010110100",  "000000101010111011",  "000000101011000011",  "000000101011001011",  "000000101011010011",  "000000101011011011",  "000000101011100011",  "000000101011101011",  "000000101011110010",  "000000101011111010",  "000000101100000010",  "000000101100001001",  "000000101100010001",  "000000101100011001",  "000000101100100000",  "000000101100101000",  "000000101100101111",  "000000101100110111",  "000000101100111110",  "000000101101000101",  "000000101101001101",  "000000101101010100",  "000000101101011100",  "000000101101100011",  "000000101101101010",  "000000101101110001",  "000000101101111001",  "000000101110000000",  "000000101110000111",  "000000101110001110",  "000000101110010101",  "000000101110011100",  "000000101110100011",  "000000101110101010",  "000000101110110001",  "000000101110111000",  "000000101110111111",  "000000101111000110",  "000000101111001101",  "000000101111010011",  "000000101111011010",  "000000101111100001",  "000000101111101000",  "000000101111101110",  "000000101111110101",  "000000101111111100",  "000000110000000010",  "000000110000001001",  "000000110000001111",  "000000110000010110",  "000000110000011100",  "000000110000100011",  "000000110000101001",  "000000110000101111",  "000000110000110110",  "000000110000111100",  "000000110001000010",  "000000110001001001",  "000000110001001111",  "000000110001010101",  "000000110001011011",  "000000110001100001",  "000000110001100111",  "000000110001101101",  "000000110001110011",  "000000110001111001",  "000000110001111111",  "000000110010000101",  "000000110010001011",  "000000110010010001",  "000000110010010111",  "000000110010011100",  "000000110010100010",  "000000110010101000",  "000000110010101110",  "000000110010110011",  "000000110010111001",  "000000110010111111",  "000000110011000100",  "000000110011001010",  "000000110011001111",  "000000110011010101",  "000000110011011010",  "000000110011011111",  "000000110011100101",  "000000110011101010",  "000000110011101111",  "000000110011110101",  "000000110011111010",  "000000110011111111",  "000000110100000100",  "000000110100001001",  "000000110100001110",  "000000110100010011",  "000000110100011001",  "000000110100011110",  "000000110100100010",  "000000110100100111",  "000000110100101100",  "000000110100110001",  "000000110100110110",  "000000110100111011",  "000000110101000000",  "000000110101000100",  "000000110101001001",  "000000110101001110",  "000000110101010010",  "000000110101010111",  "000000110101011011",  "000000110101100000",  "000000110101100100",  "000000110101101001",  "000000110101101101",  "000000110101110010",  "000000110101110110",  "000000110101111010",  "000000110101111111",  "000000110110000011",  "000000110110000111",  "000000110110001011",  "000000110110001111",  "000000110110010100",  "000000110110011000",  "000000110110011100",  "000000110110100000",  "000000110110100100",  "000000110110101000",  "000000110110101011",  "000000110110101111",  "000000110110110011",  "000000110110110111",  "000000110110111011",  "000000110110111111",  "000000110111000010",  "000000110111000110",  "000000110111001001",  "000000110111001101",  "000000110111010001",  "000000110111010100",  "000000110111011000",  "000000110111011011",  "000000110111011111",  "000000110111100010",  "000000110111100101",  "000000110111101001",  "000000110111101100",  "000000110111101111",  "000000110111110010",  "000000110111110110",  "000000110111111001",  "000000110111111100",  "000000110111111111",  "000000111000000010",  "000000111000000101",  "000000111000001000",  "000000111000001011",  "000000111000001110",  "000000111000010001",  "000000111000010011",  "000000111000010110",  "000000111000011001",  "000000111000011100",  "000000111000011110",  "000000111000100001",  "000000111000100100",  "000000111000100110",  "000000111000101001",  "000000111000101011",  "000000111000101110",  "000000111000110000",  "000000111000110011",  "000000111000110101",  "000000111000110111",  "000000111000111010",  "000000111000111100",  "000000111000111110",  "000000111001000000",  "000000111001000011",  "000000111001000101",  "000000111001000111",  "000000111001001001",  "000000111001001011",  "000000111001001101",  "000000111001001111",  "000000111001010001",  "000000111001010011",  "000000111001010100",  "000000111001010110",  "000000111001011000",  "000000111001011010",  "000000111001011011",  "000000111001011101",  "000000111001011111",  "000000111001100000",  "000000111001100010",  "000000111001100011",  "000000111001100101",  "000000111001100110",  "000000111001101000",  "000000111001101001",  "000000111001101010",  "000000111001101100",  "000000111001101101",  "000000111001101110",  "000000111001110000",  "000000111001110001",  "000000111001110010",  "000000111001110011",  "000000111001110100",  "000000111001110101",  "000000111001110110",  "000000111001110111",  "000000111001111000",  "000000111001111001",  "000000111001111010",  "000000111001111011",  "000000111001111011",  "000000111001111100",  "000000111001111101",  "000000111001111101",  "000000111001111110",  "000000111001111111",  "000000111001111111",  "000000111010000000",  "000000111010000000",  "000000111010000001",  "000000111010000001",  "000000111010000010",  "000000111010000010",  "000000111010000010",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000100",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000011",  "000000111010000010",  "000000111010000010",  "000000111010000010",  "000000111010000001",  "000000111010000001",  "000000111010000001",  "000000111010000000",  "000000111010000000",  "000000111001111111",  "000000111001111110",  "000000111001111110",  "000000111001111101",  "000000111001111101",  "000000111001111100",  "000000111001111011",  "000000111001111010",  "000000111001111001",  "000000111001111001",  "000000111001111000",  "000000111001110111",  "000000111001110110",  "000000111001110101",  "000000111001110100",  "000000111001110011",  "000000111001110010",  "000000111001110000",  "000000111001101111",  "000000111001101110",  "000000111001101101",  "000000111001101100",  "000000111001101010",  "000000111001101001",  "000000111001101000",  "000000111001100110",  "000000111001100101",  "000000111001100011",  "000000111001100010",  "000000111001100000",  "000000111001011111",  "000000111001011101",  "000000111001011011",  "000000111001011010",  "000000111001011000",  "000000111001010110",  "000000111001010100",  "000000111001010010",  "000000111001010001",  "000000111001001111",  "000000111001001101",  "000000111001001011",  "000000111001001001",  "000000111001000111",  "000000111001000101",  "000000111001000011",  "000000111001000001",  "000000111000111110",  "000000111000111100",  "000000111000111010",  "000000111000111000",  "000000111000110101",  "000000111000110011",  "000000111000110001",  "000000111000101110",  "000000111000101100",  "000000111000101001",  "000000111000100111",  "000000111000100100",  "000000111000100010",  "000000111000011111",  "000000111000011101",  "000000111000011010",  "000000111000010111",  "000000111000010101",  "000000111000010010",  "000000111000001111",  "000000111000001100",  "000000111000001001",  "000000111000000110",  "000000111000000011",  "000000111000000001",  "000000110111111110",  "000000110111111011",  "000000110111110111",  "000000110111110100",  "000000110111110001",  "000000110111101110",  "000000110111101011",  "000000110111101000",  "000000110111100100",  "000000110111100001",  "000000110111011110",  "000000110111011010",  "000000110111010111",  "000000110111010100",  "000000110111010000",  "000000110111001101",  "000000110111001001",  "000000110111000110",  "000000110111000010",  "000000110110111111",  "000000110110111011",  "000000110110110111",  "000000110110110100",  "000000110110110000",  "000000110110101100",  "000000110110101000",  "000000110110100100",  "000000110110100001",  "000000110110011101",  "000000110110011001",  "000000110110010101",  "000000110110010001",  "000000110110001101",  "000000110110001001",  "000000110110000101",  "000000110110000001",  "000000110101111100",  "000000110101111000",  "000000110101110100",  "000000110101110000",  "000000110101101100",  "000000110101100111",  "000000110101100011",  "000000110101011111",  "000000110101011010",  "000000110101010110",  "000000110101010001",  "000000110101001101",  "000000110101001000",  "000000110101000100",  "000000110100111111",  "000000110100111011",  "000000110100110110",  "000000110100110001",  "000000110100101101",  "000000110100101000",  "000000110100100011",  "000000110100011110",  "000000110100011010",  "000000110100010101",  "000000110100010000",  "000000110100001011",  "000000110100000110",  "000000110100000001",  "000000110011111100",  "000000110011110111",  "000000110011110010",  "000000110011101101",  "000000110011101000",  "000000110011100011",  "000000110011011101",  "000000110011011000",  "000000110011010011",  "000000110011001110",  "000000110011001000",  "000000110011000011",  "000000110010111110",  "000000110010111000",  "000000110010110011",  "000000110010101110",  "000000110010101000",  "000000110010100011",  "000000110010011101",  "000000110010011000",  "000000110010010010",  "000000110010001100",  "000000110010000111",  "000000110010000001",  "000000110001111011",  "000000110001110110",  "000000110001110000",  "000000110001101010",  "000000110001100100",  "000000110001011111",  "000000110001011001",  "000000110001010011",  "000000110001001101",  "000000110001000111",  "000000110001000001",  "000000110000111011",  "000000110000110101",  "000000110000101111",  "000000110000101001",  "000000110000100011",  "000000110000011101",  "000000110000010111",  "000000110000010000",  "000000110000001010",  "000000110000000100",  "000000101111111110",  "000000101111110111",  "000000101111110001",  "000000101111101011",  "000000101111100100",  "000000101111011110",  "000000101111011000",  "000000101111010001",  "000000101111001011",  "000000101111000100",  "000000101110111110",  "000000101110110111",  "000000101110110000",  "000000101110101010",  "000000101110100011",  "000000101110011101",  "000000101110010110",  "000000101110001111",  "000000101110001000",  "000000101110000010",  "000000101101111011",  "000000101101110100",  "000000101101101101",  "000000101101100110",  "000000101101100000",  "000000101101011001",  "000000101101010010",  "000000101101001011",  "000000101101000100",  "000000101100111101",  "000000101100110110",  "000000101100101111",  "000000101100101000",  "000000101100100000",  "000000101100011001",  "000000101100010010",  "000000101100001011",  "000000101100000100",  "000000101011111101",  "000000101011110101",  "000000101011101110",  "000000101011100111",  "000000101011011111",  "000000101011011000",  "000000101011010001",  "000000101011001001",  "000000101011000010",  "000000101010111010",  "000000101010110011",  "000000101010101011",  "000000101010100100",  "000000101010011100",  "000000101010010101",  "000000101010001101",  "000000101010000110",  "000000101001111110",  "000000101001110110",  "000000101001101111",  "000000101001100111",  "000000101001011111",  "000000101001011000",  "000000101001010000",  "000000101001001000",  "000000101001000000",  "000000101000111000",  "000000101000110001",  "000000101000101001",  "000000101000100001",  "000000101000011001",  "000000101000010001",  "000000101000001001",  "000000101000000001",  "000000100111111001",  "000000100111110001",  "000000100111101001",  "000000100111100001",  "000000100111011001",  "000000100111010001",  "000000100111001001",  "000000100111000001",  "000000100110111000",  "000000100110110000",  "000000100110101000",  "000000100110100000",  "000000100110010111",  "000000100110001111",  "000000100110000111",  "000000100101111111",  "000000100101110110",  "000000100101101110",  "000000100101100110",  "000000100101011101",  "000000100101010101",  "000000100101001100",  "000000100101000100",  "000000100100111011",  "000000100100110011",  "000000100100101010",  "000000100100100010",  "000000100100011001",  "000000100100010001",  "000000100100001000",  "000000100100000000",  "000000100011110111",  "000000100011101110",  "000000100011100110",  "000000100011011101",  "000000100011010100",  "000000100011001100",  "000000100011000011",  "000000100010111010",  "000000100010110001",  "000000100010101001",  "000000100010100000",  "000000100010010111",  "000000100010001110",  "000000100010000101",  "000000100001111101",  "000000100001110100",  "000000100001101011",  "000000100001100010",  "000000100001011001",  "000000100001010000",  "000000100001000111",  "000000100000111110",  "000000100000110101",  "000000100000101100",  "000000100000100011",  "000000100000011010",  "000000100000010001",  "000000100000001000",  "000000011111111111",  "000000011111110101",  "000000011111101100",  "000000011111100011",  "000000011111011010",  "000000011111010001",  "000000011111001000",  "000000011110111110",  "000000011110110101",  "000000011110101100",  "000000011110100011",  "000000011110011001",  "000000011110010000",  "000000011110000111",  "000000011101111110",  "000000011101110100",  "000000011101101011",  "000000011101100001",  "000000011101011000",  "000000011101001111",  "000000011101000101",  "000000011100111100",  "000000011100110010",  "000000011100101001",  "000000011100100000",  "000000011100010110",  "000000011100001101",  "000000011100000011",  "000000011011111010",  "000000011011110000",  "000000011011100110",  "000000011011011101",  "000000011011010011",  "000000011011001010",  "000000011011000000",  "000000011010110111",  "000000011010101101",  "000000011010100011",  "000000011010011010",  "000000011010010000",  "000000011010000110",  "000000011001111101",  "000000011001110011",  "000000011001101001",  "000000011001100000",  "000000011001010110",  "000000011001001100",  "000000011001000010",  "000000011000111001",  "000000011000101111",  "000000011000100101",  "000000011000011011",  "000000011000010001",  "000000011000001000",  "000000010111111110",  "000000010111110100",  "000000010111101010",  "000000010111100000",  "000000010111010110",  "000000010111001100",  "000000010111000010",  "000000010110111001",  "000000010110101111",  "000000010110100101",  "000000010110011011",  "000000010110010001",  "000000010110000111",  "000000010101111101",  "000000010101110011",  "000000010101101001",  "000000010101011111",  "000000010101010101",  "000000010101001011",  "000000010101000001",  "000000010100110111",  "000000010100101101",  "000000010100100011",  "000000010100011001",  "000000010100001111",  "000000010100000100",  "000000010011111010",  "000000010011110000",  "000000010011100110",  "000000010011011100",  "000000010011010010",  "000000010011001000",  "000000010010111110",  "000000010010110100",  "000000010010101001",  "000000010010011111",  "000000010010010101",  "000000010010001011",  "000000010010000001",  "000000010001110111",  "000000010001101100",  "000000010001100010",  "000000010001011000",  "000000010001001110",  "000000010001000011",  "000000010000111001",  "000000010000101111",  "000000010000100101",  "000000010000011011",  "000000010000010000",  "000000010000000110",  "000000001111111100",  "000000001111110001",  "000000001111100111",  "000000001111011101",  "000000001111010011",  "000000001111001000",  "000000001110111110",  "000000001110110100",  "000000001110101001",  "000000001110011111",  "000000001110010101",  "000000001110001010",  "000000001110000000",  "000000001101110110",  "000000001101101011",  "000000001101100001",  "000000001101010111",  "000000001101001100",  "000000001101000010",  "000000001100111000",  "000000001100101101",  "000000001100100011",  "000000001100011000",  "000000001100001110",  "000000001100000100",  "000000001011111001",  "000000001011101111",  "000000001011100101",  "000000001011011010",  "000000001011010000",  "000000001011000101",  "000000001010111011",  "000000001010110001",  "000000001010100110",  "000000001010011100",  "000000001010010001",  "000000001010000111",  "000000001001111100",  "000000001001110010",  "000000001001101000",  "000000001001011101",  "000000001001010011",  "000000001001001000",  "000000001000111110",  "000000001000110011",  "000000001000101001",  "000000001000011111",  "000000001000010100",  "000000001000001010",  "000000000111111111",  "000000000111110101",  "000000000111101010",  "000000000111100000",  "000000000111010101",  "000000000111001011",  "000000000111000000",  "000000000110110110",  "000000000110101100",  "000000000110100001",  "000000000110010111",  "000000000110001100",  "000000000110000010",  "000000000101110111",  "000000000101101101",  "000000000101100010",  "000000000101011000",  "000000000101001110",  "000000000101000011",  "000000000100111001",  "000000000100101110",  "000000000100100100",  "000000000100011001",  "000000000100001111",  "000000000100000100",  "000000000011111010",  "000000000011110000",  "000000000011100101",  "000000000011011011",  "000000000011010000",  "000000000011000110",  "000000000010111011",  "000000000010110001",  "000000000010100110",  "000000000010011100",  "000000000010010010",  "000000000010000111",  "000000000001111101",  "000000000001110010",  "000000000001101000",  "000000000001011110",  "000000000001010011",  "000000000001001001",  "000000000000111110",  "000000000000110100",  "000000000000101010",  "000000000000011111",  "000000000000010101",  "000000000000001010"),("000000000000000000",  "111111111111110110",  "111111111111101011",  "111111111111100001",  "111111111111010111",  "111111111111001100",  "111111111111000010",  "111111111110110111",  "111111111110101101",  "111111111110100011",  "111111111110011000",  "111111111110001110",  "111111111110000100",  "111111111101111001",  "111111111101101111",  "111111111101100101",  "111111111101011010",  "111111111101010000",  "111111111101000110",  "111111111100111100",  "111111111100110001",  "111111111100100111",  "111111111100011101",  "111111111100010010",  "111111111100001000",  "111111111011111110",  "111111111011110100",  "111111111011101001",  "111111111011011111",  "111111111011010101",  "111111111011001011",  "111111111011000000",  "111111111010110110",  "111111111010101100",  "111111111010100010",  "111111111010011000",  "111111111010001101",  "111111111010000011",  "111111111001111001",  "111111111001101111",  "111111111001100101",  "111111111001011011",  "111111111001010000",  "111111111001000110",  "111111111000111100",  "111111111000110010",  "111111111000101000",  "111111111000011110",  "111111111000010100",  "111111111000001010",  "111111111000000000",  "111111110111110110",  "111111110111101011",  "111111110111100001",  "111111110111010111",  "111111110111001101",  "111111110111000011",  "111111110110111001",  "111111110110101111",  "111111110110100101",  "111111110110011011",  "111111110110010001",  "111111110110000111",  "111111110101111101",  "111111110101110011",  "111111110101101001",  "111111110101100000",  "111111110101010110",  "111111110101001100",  "111111110101000010",  "111111110100111000",  "111111110100101110",  "111111110100100100",  "111111110100011010",  "111111110100010000",  "111111110100000111",  "111111110011111101",  "111111110011110011",  "111111110011101001",  "111111110011011111",  "111111110011010110",  "111111110011001100",  "111111110011000010",  "111111110010111000",  "111111110010101110",  "111111110010100101",  "111111110010011011",  "111111110010010001",  "111111110010001000",  "111111110001111110",  "111111110001110100",  "111111110001101011",  "111111110001100001",  "111111110001010111",  "111111110001001110",  "111111110001000100",  "111111110000111010",  "111111110000110001",  "111111110000100111",  "111111110000011110",  "111111110000010100",  "111111110000001011",  "111111110000000001",  "111111101111111000",  "111111101111101110",  "111111101111100101",  "111111101111011011",  "111111101111010010",  "111111101111001000",  "111111101110111111",  "111111101110110101",  "111111101110101100",  "111111101110100011",  "111111101110011001",  "111111101110010000",  "111111101110000111",  "111111101101111101",  "111111101101110100",  "111111101101101011",  "111111101101100001",  "111111101101011000",  "111111101101001111",  "111111101101000110",  "111111101100111100",  "111111101100110011",  "111111101100101010",  "111111101100100001",  "111111101100011000",  "111111101100001110",  "111111101100000101",  "111111101011111100",  "111111101011110011",  "111111101011101010",  "111111101011100001",  "111111101011011000",  "111111101011001111",  "111111101011000110",  "111111101010111101",  "111111101010110100",  "111111101010101011",  "111111101010100010",  "111111101010011001",  "111111101010010000",  "111111101010000111",  "111111101001111110",  "111111101001110101",  "111111101001101100",  "111111101001100011",  "111111101001011011",  "111111101001010010",  "111111101001001001",  "111111101001000000",  "111111101000110111",  "111111101000101111",  "111111101000100110",  "111111101000011101",  "111111101000010101",  "111111101000001100",  "111111101000000011",  "111111100111111011",  "111111100111110010",  "111111100111101001",  "111111100111100001",  "111111100111011000",  "111111100111010000",  "111111100111000111",  "111111100110111110",  "111111100110110110",  "111111100110101101",  "111111100110100101",  "111111100110011101",  "111111100110010100",  "111111100110001100",  "111111100110000011",  "111111100101111011",  "111111100101110011",  "111111100101101010",  "111111100101100010",  "111111100101011010",  "111111100101010001",  "111111100101001001",  "111111100101000001",  "111111100100111001",  "111111100100110000",  "111111100100101000",  "111111100100100000",  "111111100100011000",  "111111100100010000",  "111111100100001000",  "111111100100000000",  "111111100011111000",  "111111100011101111",  "111111100011100111",  "111111100011011111",  "111111100011010111",  "111111100011001111",  "111111100011001000",  "111111100011000000",  "111111100010111000",  "111111100010110000",  "111111100010101000",  "111111100010100000",  "111111100010011000",  "111111100010010000",  "111111100010001001",  "111111100010000001",  "111111100001111001",  "111111100001110001",  "111111100001101010",  "111111100001100010",  "111111100001011010",  "111111100001010011",  "111111100001001011",  "111111100001000100",  "111111100000111100",  "111111100000110100",  "111111100000101101",  "111111100000100101",  "111111100000011110",  "111111100000010110",  "111111100000001111",  "111111100000001000",  "111111100000000000",  "111111011111111001",  "111111011111110001",  "111111011111101010",  "111111011111100011",  "111111011111011100",  "111111011111010100",  "111111011111001101",  "111111011111000110",  "111111011110111111",  "111111011110110111",  "111111011110110000",  "111111011110101001",  "111111011110100010",  "111111011110011011",  "111111011110010100",  "111111011110001101",  "111111011110000110",  "111111011101111111",  "111111011101111000",  "111111011101110001",  "111111011101101010",  "111111011101100011",  "111111011101011100",  "111111011101010101",  "111111011101001111",  "111111011101001000",  "111111011101000001",  "111111011100111010",  "111111011100110011",  "111111011100101101",  "111111011100100110",  "111111011100011111",  "111111011100011001",  "111111011100010010",  "111111011100001100",  "111111011100000101",  "111111011011111110",  "111111011011111000",  "111111011011110001",  "111111011011101011",  "111111011011100100",  "111111011011011110",  "111111011011011000",  "111111011011010001",  "111111011011001011",  "111111011011000101",  "111111011010111110",  "111111011010111000",  "111111011010110010",  "111111011010101100",  "111111011010100101",  "111111011010011111",  "111111011010011001",  "111111011010010011",  "111111011010001101",  "111111011010000111",  "111111011010000001",  "111111011001111011",  "111111011001110101",  "111111011001101111",  "111111011001101001",  "111111011001100011",  "111111011001011101",  "111111011001010111",  "111111011001010001",  "111111011001001011",  "111111011001000101",  "111111011001000000",  "111111011000111010",  "111111011000110100",  "111111011000101110",  "111111011000101001",  "111111011000100011",  "111111011000011110",  "111111011000011000",  "111111011000010010",  "111111011000001101",  "111111011000000111",  "111111011000000010",  "111111010111111100",  "111111010111110111",  "111111010111110010",  "111111010111101100",  "111111010111100111",  "111111010111100001",  "111111010111011100",  "111111010111010111",  "111111010111010010",  "111111010111001100",  "111111010111000111",  "111111010111000010",  "111111010110111101",  "111111010110111000",  "111111010110110011",  "111111010110101110",  "111111010110101000",  "111111010110100011",  "111111010110011110",  "111111010110011010",  "111111010110010101",  "111111010110010000",  "111111010110001011",  "111111010110000110",  "111111010110000001",  "111111010101111100",  "111111010101111000",  "111111010101110011",  "111111010101101110",  "111111010101101001",  "111111010101100101",  "111111010101100000",  "111111010101011011",  "111111010101010111",  "111111010101010010",  "111111010101001110",  "111111010101001001",  "111111010101000101",  "111111010101000000",  "111111010100111100",  "111111010100111000",  "111111010100110011",  "111111010100101111",  "111111010100101011",  "111111010100100110",  "111111010100100010",  "111111010100011110",  "111111010100011010",  "111111010100010101",  "111111010100010001",  "111111010100001101",  "111111010100001001",  "111111010100000101",  "111111010100000001",  "111111010011111101",  "111111010011111001",  "111111010011110101",  "111111010011110001",  "111111010011101101",  "111111010011101001",  "111111010011100110",  "111111010011100010",  "111111010011011110",  "111111010011011010",  "111111010011010111",  "111111010011010011",  "111111010011001111",  "111111010011001100",  "111111010011001000",  "111111010011000100",  "111111010011000001",  "111111010010111101",  "111111010010111010",  "111111010010110110",  "111111010010110011",  "111111010010110000",  "111111010010101100",  "111111010010101001",  "111111010010100101",  "111111010010100010",  "111111010010011111",  "111111010010011100",  "111111010010011000",  "111111010010010101",  "111111010010010010",  "111111010010001111",  "111111010010001100",  "111111010010001001",  "111111010010000110",  "111111010010000011",  "111111010010000000",  "111111010001111101",  "111111010001111010",  "111111010001110111",  "111111010001110100",  "111111010001110001",  "111111010001101111",  "111111010001101100",  "111111010001101001",  "111111010001100110",  "111111010001100100",  "111111010001100001",  "111111010001011110",  "111111010001011100",  "111111010001011001",  "111111010001010111",  "111111010001010100",  "111111010001010010",  "111111010001001111",  "111111010001001101",  "111111010001001010",  "111111010001001000",  "111111010001000110",  "111111010001000011",  "111111010001000001",  "111111010000111111",  "111111010000111101",  "111111010000111010",  "111111010000111000",  "111111010000110110",  "111111010000110100",  "111111010000110010",  "111111010000110000",  "111111010000101110",  "111111010000101100",  "111111010000101010",  "111111010000101000",  "111111010000100110",  "111111010000100100",  "111111010000100010",  "111111010000100001",  "111111010000011111",  "111111010000011101",  "111111010000011011",  "111111010000011010",  "111111010000011000",  "111111010000010110",  "111111010000010101",  "111111010000010011",  "111111010000010010",  "111111010000010000",  "111111010000001111",  "111111010000001101",  "111111010000001100",  "111111010000001010",  "111111010000001001",  "111111010000001000",  "111111010000000110",  "111111010000000101",  "111111010000000100",  "111111010000000011",  "111111010000000001",  "111111010000000000",  "111111001111111111",  "111111001111111110",  "111111001111111101",  "111111001111111100",  "111111001111111011",  "111111001111111010",  "111111001111111001",  "111111001111111000",  "111111001111110111",  "111111001111110110",  "111111001111110101",  "111111001111110100",  "111111001111110100",  "111111001111110011",  "111111001111110010",  "111111001111110010",  "111111001111110001",  "111111001111110000",  "111111001111110000",  "111111001111101111",  "111111001111101110",  "111111001111101110",  "111111001111101101",  "111111001111101101",  "111111001111101101",  "111111001111101100",  "111111001111101100",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101010",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101011",  "111111001111101100",  "111111001111101100",  "111111001111101100",  "111111001111101101",  "111111001111101101",  "111111001111101110",  "111111001111101110",  "111111001111101111",  "111111001111101111",  "111111001111110000",  "111111001111110001",  "111111001111110001",  "111111001111110010",  "111111001111110011",  "111111001111110011",  "111111001111110100",  "111111001111110101",  "111111001111110110",  "111111001111110111",  "111111001111110111",  "111111001111111000",  "111111001111111001",  "111111001111111010",  "111111001111111011",  "111111001111111100",  "111111001111111101",  "111111001111111110",  "111111001111111111",  "111111010000000001",  "111111010000000010",  "111111010000000011",  "111111010000000100",  "111111010000000101",  "111111010000000111",  "111111010000001000",  "111111010000001001",  "111111010000001011",  "111111010000001100",  "111111010000001110",  "111111010000001111",  "111111010000010000",  "111111010000010010",  "111111010000010100",  "111111010000010101",  "111111010000010111",  "111111010000011000",  "111111010000011010",  "111111010000011100",  "111111010000011101",  "111111010000011111",  "111111010000100001",  "111111010000100011",  "111111010000100100",  "111111010000100110",  "111111010000101000",  "111111010000101010",  "111111010000101100",  "111111010000101110",  "111111010000110000",  "111111010000110010",  "111111010000110100",  "111111010000110110",  "111111010000111000",  "111111010000111010",  "111111010000111100",  "111111010000111111",  "111111010001000001",  "111111010001000011",  "111111010001000101",  "111111010001001000",  "111111010001001010",  "111111010001001100",  "111111010001001111",  "111111010001010001",  "111111010001010011",  "111111010001010110",  "111111010001011000",  "111111010001011011",  "111111010001011101",  "111111010001100000",  "111111010001100011",  "111111010001100101",  "111111010001101000",  "111111010001101011",  "111111010001101101",  "111111010001110000",  "111111010001110011",  "111111010001110101",  "111111010001111000",  "111111010001111011",  "111111010001111110",  "111111010010000001",  "111111010010000100",  "111111010010000111",  "111111010010001010",  "111111010010001101",  "111111010010010000",  "111111010010010011",  "111111010010010110",  "111111010010011001",  "111111010010011100",  "111111010010011111",  "111111010010100010",  "111111010010100110",  "111111010010101001",  "111111010010101100",  "111111010010101111",  "111111010010110011",  "111111010010110110",  "111111010010111001",  "111111010010111101",  "111111010011000000",  "111111010011000100",  "111111010011000111",  "111111010011001011",  "111111010011001110",  "111111010011010010",  "111111010011010101",  "111111010011011001",  "111111010011011100",  "111111010011100000",  "111111010011100100",  "111111010011100111",  "111111010011101011",  "111111010011101111",  "111111010011110011",  "111111010011110110",  "111111010011111010",  "111111010011111110",  "111111010100000010",  "111111010100000110",  "111111010100001010",  "111111010100001110",  "111111010100010010",  "111111010100010110",  "111111010100011010",  "111111010100011110",  "111111010100100010",  "111111010100100110",  "111111010100101010",  "111111010100101110",  "111111010100110011",  "111111010100110111",  "111111010100111011",  "111111010100111111",  "111111010101000011",  "111111010101001000",  "111111010101001100",  "111111010101010000",  "111111010101010101",  "111111010101011001",  "111111010101011110",  "111111010101100010",  "111111010101100111",  "111111010101101011",  "111111010101110000",  "111111010101110100",  "111111010101111001",  "111111010101111101",  "111111010110000010",  "111111010110000110",  "111111010110001011",  "111111010110010000",  "111111010110010101",  "111111010110011001",  "111111010110011110",  "111111010110100011",  "111111010110101000",  "111111010110101100",  "111111010110110001",  "111111010110110110",  "111111010110111011",  "111111010111000000",  "111111010111000101",  "111111010111001010",  "111111010111001111",  "111111010111010100",  "111111010111011001",  "111111010111011110",  "111111010111100011",  "111111010111101000",  "111111010111101101",  "111111010111110010",  "111111010111110111",  "111111010111111101",  "111111011000000010",  "111111011000000111",  "111111011000001100",  "111111011000010010",  "111111011000010111",  "111111011000011100",  "111111011000100010",  "111111011000100111",  "111111011000101100",  "111111011000110010",  "111111011000110111",  "111111011000111101",  "111111011001000010",  "111111011001001000",  "111111011001001101",  "111111011001010011",  "111111011001011000",  "111111011001011110",  "111111011001100011",  "111111011001101001",  "111111011001101111",  "111111011001110100",  "111111011001111010",  "111111011010000000",  "111111011010000101",  "111111011010001011",  "111111011010010001",  "111111011010010111",  "111111011010011101",  "111111011010100010",  "111111011010101000",  "111111011010101110",  "111111011010110100",  "111111011010111010",  "111111011011000000",  "111111011011000110",  "111111011011001100",  "111111011011010010",  "111111011011011000",  "111111011011011110",  "111111011011100100",  "111111011011101010",  "111111011011110000",  "111111011011110110",  "111111011011111100",  "111111011100000011",  "111111011100001001",  "111111011100001111",  "111111011100010101",  "111111011100011011",  "111111011100100010",  "111111011100101000",  "111111011100101110",  "111111011100110100",  "111111011100111011",  "111111011101000001",  "111111011101001000",  "111111011101001110",  "111111011101010100",  "111111011101011011",  "111111011101100001",  "111111011101101000",  "111111011101101110",  "111111011101110101",  "111111011101111011",  "111111011110000010",  "111111011110001000",  "111111011110001111",  "111111011110010101",  "111111011110011100",  "111111011110100011",  "111111011110101001",  "111111011110110000",  "111111011110110111",  "111111011110111101",  "111111011111000100",  "111111011111001011",  "111111011111010001",  "111111011111011000",  "111111011111011111",  "111111011111100110",  "111111011111101101",  "111111011111110011",  "111111011111111010",  "111111100000000001",  "111111100000001000",  "111111100000001111",  "111111100000010110",  "111111100000011101",  "111111100000100100",  "111111100000101011",  "111111100000110010",  "111111100000111001",  "111111100001000000",  "111111100001000111",  "111111100001001110",  "111111100001010101",  "111111100001011100",  "111111100001100011",  "111111100001101010",  "111111100001110001",  "111111100001111000",  "111111100010000000",  "111111100010000111",  "111111100010001110",  "111111100010010101",  "111111100010011100",  "111111100010100100",  "111111100010101011",  "111111100010110010",  "111111100010111001",  "111111100011000001",  "111111100011001000",  "111111100011001111",  "111111100011010111",  "111111100011011110",  "111111100011100101",  "111111100011101101",  "111111100011110100",  "111111100011111100",  "111111100100000011",  "111111100100001011",  "111111100100010010",  "111111100100011010",  "111111100100100001",  "111111100100101000",  "111111100100110000",  "111111100100111000",  "111111100100111111",  "111111100101000111",  "111111100101001110",  "111111100101010110",  "111111100101011101",  "111111100101100101",  "111111100101101101",  "111111100101110100",  "111111100101111100",  "111111100110000100",  "111111100110001011",  "111111100110010011",  "111111100110011011",  "111111100110100010",  "111111100110101010",  "111111100110110010",  "111111100110111010",  "111111100111000001",  "111111100111001001",  "111111100111010001",  "111111100111011001",  "111111100111100001",  "111111100111101000",  "111111100111110000",  "111111100111111000",  "111111101000000000",  "111111101000001000",  "111111101000010000",  "111111101000011000",  "111111101000011111",  "111111101000100111",  "111111101000101111",  "111111101000110111",  "111111101000111111",  "111111101001000111",  "111111101001001111",  "111111101001010111",  "111111101001011111",  "111111101001100111",  "111111101001101111",  "111111101001110111",  "111111101001111111",  "111111101010000111",  "111111101010001111",  "111111101010010111",  "111111101010011111",  "111111101010101000",  "111111101010110000",  "111111101010111000",  "111111101011000000",  "111111101011001000",  "111111101011010000",  "111111101011011000",  "111111101011100000",  "111111101011101001",  "111111101011110001",  "111111101011111001",  "111111101100000001",  "111111101100001001",  "111111101100010010",  "111111101100011010",  "111111101100100010",  "111111101100101010",  "111111101100110011",  "111111101100111011",  "111111101101000011",  "111111101101001011",  "111111101101010100",  "111111101101011100",  "111111101101100100",  "111111101101101101",  "111111101101110101",  "111111101101111101",  "111111101110000110",  "111111101110001110",  "111111101110010110",  "111111101110011111",  "111111101110100111",  "111111101110101111",  "111111101110111000",  "111111101111000000",  "111111101111001001",  "111111101111010001",  "111111101111011001",  "111111101111100010",  "111111101111101010",  "111111101111110011",  "111111101111111011",  "111111110000000011",  "111111110000001100",  "111111110000010100",  "111111110000011101",  "111111110000100101",  "111111110000101110",  "111111110000110110",  "111111110000111111",  "111111110001000111",  "111111110001010000",  "111111110001011000",  "111111110001100001",  "111111110001101001",  "111111110001110010",  "111111110001111010",  "111111110010000011",  "111111110010001011",  "111111110010010100",  "111111110010011101",  "111111110010100101",  "111111110010101110",  "111111110010110110",  "111111110010111111",  "111111110011000111",  "111111110011010000",  "111111110011011001",  "111111110011100001",  "111111110011101010",  "111111110011110010",  "111111110011111011",  "111111110100000100",  "111111110100001100",  "111111110100010101",  "111111110100011101",  "111111110100100110",  "111111110100101111",  "111111110100110111",  "111111110101000000",  "111111110101001001",  "111111110101010001",  "111111110101011010",  "111111110101100010",  "111111110101101011",  "111111110101110100",  "111111110101111100",  "111111110110000101",  "111111110110001110",  "111111110110010110",  "111111110110011111",  "111111110110101000",  "111111110110110000",  "111111110110111001",  "111111110111000010",  "111111110111001010",  "111111110111010011",  "111111110111011100",  "111111110111100101",  "111111110111101101",  "111111110111110110",  "111111110111111111",  "111111111000000111",  "111111111000010000",  "111111111000011001",  "111111111000100001",  "111111111000101010",  "111111111000110011",  "111111111000111100",  "111111111001000100",  "111111111001001101",  "111111111001010110",  "111111111001011110",  "111111111001100111",  "111111111001110000",  "111111111001111001",  "111111111010000001",  "111111111010001010",  "111111111010010011",  "111111111010011011",  "111111111010100100",  "111111111010101101",  "111111111010110110",  "111111111010111110",  "111111111011000111",  "111111111011010000",  "111111111011011000",  "111111111011100001",  "111111111011101010",  "111111111011110011",  "111111111011111011",  "111111111100000100",  "111111111100001101",  "111111111100010101",  "111111111100011110",  "111111111100100111",  "111111111100110000",  "111111111100111000",  "111111111101000001",  "111111111101001010",  "111111111101010010",  "111111111101011011",  "111111111101100100",  "111111111101101100",  "111111111101110101",  "111111111101111110",  "111111111110000111",  "111111111110001111",  "111111111110011000",  "111111111110100001",  "111111111110101001",  "111111111110110010",  "111111111110111011",  "111111111111000011",  "111111111111001100",  "111111111111010101",  "111111111111011101",  "111111111111100110",  "111111111111101111",  "111111111111110111"),("000000000000000000",  "000000000000001001",  "000000000000010001",  "000000000000011010",  "000000000000100011",  "000000000000101011",  "000000000000110100",  "000000000000111101",  "000000000001000101",  "000000000001001110",  "000000000001010110",  "000000000001011111",  "000000000001101000",  "000000000001110000",  "000000000001111001",  "000000000010000001",  "000000000010001010",  "000000000010010011",  "000000000010011011",  "000000000010100100",  "000000000010101100",  "000000000010110101",  "000000000010111110",  "000000000011000110",  "000000000011001111",  "000000000011010111",  "000000000011100000",  "000000000011101000",  "000000000011110001",  "000000000011111001",  "000000000100000010",  "000000000100001011",  "000000000100010011",  "000000000100011100",  "000000000100100100",  "000000000100101101",  "000000000100110101",  "000000000100111110",  "000000000101000110",  "000000000101001111",  "000000000101010111",  "000000000101100000",  "000000000101101000",  "000000000101110000",  "000000000101111001",  "000000000110000001",  "000000000110001010",  "000000000110010010",  "000000000110011011",  "000000000110100011",  "000000000110101011",  "000000000110110100",  "000000000110111100",  "000000000111000101",  "000000000111001101",  "000000000111010101",  "000000000111011110",  "000000000111100110",  "000000000111101110",  "000000000111110111",  "000000000111111111",  "000000001000000111",  "000000001000010000",  "000000001000011000",  "000000001000100000",  "000000001000101001",  "000000001000110001",  "000000001000111001",  "000000001001000010",  "000000001001001010",  "000000001001010010",  "000000001001011010",  "000000001001100011",  "000000001001101011",  "000000001001110011",  "000000001001111011",  "000000001010000011",  "000000001010001100",  "000000001010010100",  "000000001010011100",  "000000001010100100",  "000000001010101100",  "000000001010110100",  "000000001010111101",  "000000001011000101",  "000000001011001101",  "000000001011010101",  "000000001011011101",  "000000001011100101",  "000000001011101101",  "000000001011110101",  "000000001011111101",  "000000001100000101",  "000000001100001101",  "000000001100010101",  "000000001100011101",  "000000001100100110",  "000000001100101110",  "000000001100110101",  "000000001100111101",  "000000001101000101",  "000000001101001101",  "000000001101010101",  "000000001101011101",  "000000001101100101",  "000000001101101101",  "000000001101110101",  "000000001101111101",  "000000001110000101",  "000000001110001101",  "000000001110010101",  "000000001110011100",  "000000001110100100",  "000000001110101100",  "000000001110110100",  "000000001110111100",  "000000001111000011",  "000000001111001011",  "000000001111010011",  "000000001111011011",  "000000001111100010",  "000000001111101010",  "000000001111110010",  "000000001111111010",  "000000010000000001",  "000000010000001001",  "000000010000010001",  "000000010000011000",  "000000010000100000",  "000000010000101000",  "000000010000101111",  "000000010000110111",  "000000010000111110",  "000000010001000110",  "000000010001001110",  "000000010001010101",  "000000010001011101",  "000000010001100100",  "000000010001101100",  "000000010001110011",  "000000010001111011",  "000000010010000010",  "000000010010001010",  "000000010010010001",  "000000010010011000",  "000000010010100000",  "000000010010100111",  "000000010010101111",  "000000010010110110",  "000000010010111101",  "000000010011000101",  "000000010011001100",  "000000010011010011",  "000000010011011011",  "000000010011100010",  "000000010011101001",  "000000010011110001",  "000000010011111000",  "000000010011111111",  "000000010100000110",  "000000010100001101",  "000000010100010101",  "000000010100011100",  "000000010100100011",  "000000010100101010",  "000000010100110001",  "000000010100111000",  "000000010100111111",  "000000010101000111",  "000000010101001110",  "000000010101010101",  "000000010101011100",  "000000010101100011",  "000000010101101010",  "000000010101110001",  "000000010101111000",  "000000010101111111",  "000000010110000110",  "000000010110001100",  "000000010110010011",  "000000010110011010",  "000000010110100001",  "000000010110101000",  "000000010110101111",  "000000010110110110",  "000000010110111101",  "000000010111000011",  "000000010111001010",  "000000010111010001",  "000000010111011000",  "000000010111011110",  "000000010111100101",  "000000010111101100",  "000000010111110010",  "000000010111111001",  "000000011000000000",  "000000011000000110",  "000000011000001101",  "000000011000010100",  "000000011000011010",  "000000011000100001",  "000000011000100111",  "000000011000101110",  "000000011000110100",  "000000011000111011",  "000000011001000001",  "000000011001001000",  "000000011001001110",  "000000011001010101",  "000000011001011011",  "000000011001100010",  "000000011001101000",  "000000011001101110",  "000000011001110101",  "000000011001111011",  "000000011010000001",  "000000011010001000",  "000000011010001110",  "000000011010010100",  "000000011010011010",  "000000011010100000",  "000000011010100111",  "000000011010101101",  "000000011010110011",  "000000011010111001",  "000000011010111111",  "000000011011000101",  "000000011011001011",  "000000011011010010",  "000000011011011000",  "000000011011011110",  "000000011011100100",  "000000011011101010",  "000000011011110000",  "000000011011110110",  "000000011011111011",  "000000011100000001",  "000000011100000111",  "000000011100001101",  "000000011100010011",  "000000011100011001",  "000000011100011111",  "000000011100100100",  "000000011100101010",  "000000011100110000",  "000000011100110110",  "000000011100111011",  "000000011101000001",  "000000011101000111",  "000000011101001101",  "000000011101010010",  "000000011101011000",  "000000011101011101",  "000000011101100011",  "000000011101101001",  "000000011101101110",  "000000011101110100",  "000000011101111001",  "000000011101111111",  "000000011110000100",  "000000011110001010",  "000000011110001111",  "000000011110010100",  "000000011110011010",  "000000011110011111",  "000000011110100100",  "000000011110101010",  "000000011110101111",  "000000011110110100",  "000000011110111010",  "000000011110111111",  "000000011111000100",  "000000011111001001",  "000000011111001111",  "000000011111010100",  "000000011111011001",  "000000011111011110",  "000000011111100011",  "000000011111101000",  "000000011111101101",  "000000011111110010",  "000000011111110111",  "000000011111111100",  "000000100000000001",  "000000100000000110",  "000000100000001011",  "000000100000010000",  "000000100000010101",  "000000100000011010",  "000000100000011111",  "000000100000100011",  "000000100000101000",  "000000100000101101",  "000000100000110010",  "000000100000110110",  "000000100000111011",  "000000100001000000",  "000000100001000101",  "000000100001001001",  "000000100001001110",  "000000100001010010",  "000000100001010111",  "000000100001011100",  "000000100001100000",  "000000100001100101",  "000000100001101001",  "000000100001101110",  "000000100001110010",  "000000100001110111",  "000000100001111011",  "000000100001111111",  "000000100010000100",  "000000100010001000",  "000000100010001100",  "000000100010010001",  "000000100010010101",  "000000100010011001",  "000000100010011101",  "000000100010100010",  "000000100010100110",  "000000100010101010",  "000000100010101110",  "000000100010110010",  "000000100010110110",  "000000100010111010",  "000000100010111111",  "000000100011000011",  "000000100011000111",  "000000100011001011",  "000000100011001111",  "000000100011010010",  "000000100011010110",  "000000100011011010",  "000000100011011110",  "000000100011100010",  "000000100011100110",  "000000100011101010",  "000000100011101101",  "000000100011110001",  "000000100011110101",  "000000100011111001",  "000000100011111100",  "000000100100000000",  "000000100100000100",  "000000100100000111",  "000000100100001011",  "000000100100001110",  "000000100100010010",  "000000100100010110",  "000000100100011001",  "000000100100011101",  "000000100100100000",  "000000100100100011",  "000000100100100111",  "000000100100101010",  "000000100100101110",  "000000100100110001",  "000000100100110100",  "000000100100111000",  "000000100100111011",  "000000100100111110",  "000000100101000001",  "000000100101000100",  "000000100101001000",  "000000100101001011",  "000000100101001110",  "000000100101010001",  "000000100101010100",  "000000100101010111",  "000000100101011010",  "000000100101011101",  "000000100101100000",  "000000100101100011",  "000000100101100110",  "000000100101101001",  "000000100101101100",  "000000100101101111",  "000000100101110010",  "000000100101110101",  "000000100101110111",  "000000100101111010",  "000000100101111101",  "000000100110000000",  "000000100110000010",  "000000100110000101",  "000000100110001000",  "000000100110001010",  "000000100110001101",  "000000100110001111",  "000000100110010010",  "000000100110010101",  "000000100110010111",  "000000100110011010",  "000000100110011100",  "000000100110011110",  "000000100110100001",  "000000100110100011",  "000000100110100110",  "000000100110101000",  "000000100110101010",  "000000100110101101",  "000000100110101111",  "000000100110110001",  "000000100110110011",  "000000100110110110",  "000000100110111000",  "000000100110111010",  "000000100110111100",  "000000100110111110",  "000000100111000000",  "000000100111000010",  "000000100111000100",  "000000100111000110",  "000000100111001000",  "000000100111001010",  "000000100111001100",  "000000100111001110",  "000000100111010000",  "000000100111010010",  "000000100111010100",  "000000100111010101",  "000000100111010111",  "000000100111011001",  "000000100111011011",  "000000100111011100",  "000000100111011110",  "000000100111100000",  "000000100111100001",  "000000100111100011",  "000000100111100101",  "000000100111100110",  "000000100111101000",  "000000100111101001",  "000000100111101011",  "000000100111101100",  "000000100111101110",  "000000100111101111",  "000000100111110000",  "000000100111110010",  "000000100111110011",  "000000100111110100",  "000000100111110110",  "000000100111110111",  "000000100111111000",  "000000100111111001",  "000000100111111011",  "000000100111111100",  "000000100111111101",  "000000100111111110",  "000000100111111111",  "000000101000000000",  "000000101000000001",  "000000101000000010",  "000000101000000011",  "000000101000000100",  "000000101000000101",  "000000101000000110",  "000000101000000111",  "000000101000001000",  "000000101000001001",  "000000101000001010",  "000000101000001010",  "000000101000001011",  "000000101000001100",  "000000101000001101",  "000000101000001101",  "000000101000001110",  "000000101000001111",  "000000101000001111",  "000000101000010000",  "000000101000010001",  "000000101000010001",  "000000101000010010",  "000000101000010010",  "000000101000010011",  "000000101000010011",  "000000101000010100",  "000000101000010100",  "000000101000010100",  "000000101000010101",  "000000101000010101",  "000000101000010101",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010111",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010110",  "000000101000010101",  "000000101000010101",  "000000101000010101",  "000000101000010100",  "000000101000010100",  "000000101000010011",  "000000101000010011",  "000000101000010011",  "000000101000010010",  "000000101000010010",  "000000101000010001",  "000000101000010000",  "000000101000010000",  "000000101000001111",  "000000101000001111",  "000000101000001110",  "000000101000001101",  "000000101000001101",  "000000101000001100",  "000000101000001011",  "000000101000001010",  "000000101000001001",  "000000101000001001",  "000000101000001000",  "000000101000000111",  "000000101000000110",  "000000101000000101",  "000000101000000100",  "000000101000000011",  "000000101000000010",  "000000101000000001",  "000000101000000000",  "000000100111111111",  "000000100111111110",  "000000100111111101",  "000000100111111100",  "000000100111111011",  "000000100111111001",  "000000100111111000",  "000000100111110111",  "000000100111110110",  "000000100111110100",  "000000100111110011",  "000000100111110010",  "000000100111110000",  "000000100111101111",  "000000100111101110",  "000000100111101100",  "000000100111101011",  "000000100111101001",  "000000100111101000",  "000000100111100110",  "000000100111100101",  "000000100111100011",  "000000100111100010",  "000000100111100000",  "000000100111011110",  "000000100111011101",  "000000100111011011",  "000000100111011001",  "000000100111011000",  "000000100111010110",  "000000100111010100",  "000000100111010010",  "000000100111010001",  "000000100111001111",  "000000100111001101",  "000000100111001011",  "000000100111001001",  "000000100111000111",  "000000100111000101",  "000000100111000011",  "000000100111000001",  "000000100110111111",  "000000100110111101",  "000000100110111011",  "000000100110111001",  "000000100110110111",  "000000100110110101",  "000000100110110011",  "000000100110110000",  "000000100110101110",  "000000100110101100",  "000000100110101010",  "000000100110100111",  "000000100110100101",  "000000100110100011",  "000000100110100000",  "000000100110011110",  "000000100110011100",  "000000100110011001",  "000000100110010111",  "000000100110010100",  "000000100110010010",  "000000100110001111",  "000000100110001101",  "000000100110001010",  "000000100110001000",  "000000100110000101",  "000000100110000011",  "000000100110000000",  "000000100101111101",  "000000100101111011",  "000000100101111000",  "000000100101110101",  "000000100101110010",  "000000100101110000",  "000000100101101101",  "000000100101101010",  "000000100101100111",  "000000100101100100",  "000000100101100010",  "000000100101011111",  "000000100101011100",  "000000100101011001",  "000000100101010110",  "000000100101010011",  "000000100101010000",  "000000100101001101",  "000000100101001010",  "000000100101000111",  "000000100101000100",  "000000100101000001",  "000000100100111101",  "000000100100111010",  "000000100100110111",  "000000100100110100",  "000000100100110001",  "000000100100101110",  "000000100100101010",  "000000100100100111",  "000000100100100100",  "000000100100100000",  "000000100100011101",  "000000100100011010",  "000000100100010110",  "000000100100010011",  "000000100100001111",  "000000100100001100",  "000000100100001001",  "000000100100000101",  "000000100100000010",  "000000100011111110",  "000000100011111010",  "000000100011110111",  "000000100011110011",  "000000100011110000",  "000000100011101100",  "000000100011101000",  "000000100011100101",  "000000100011100001",  "000000100011011101",  "000000100011011010",  "000000100011010110",  "000000100011010010",  "000000100011001110",  "000000100011001011",  "000000100011000111",  "000000100011000011",  "000000100010111111",  "000000100010111011",  "000000100010110111",  "000000100010110011",  "000000100010101111",  "000000100010101011",  "000000100010100111",  "000000100010100011",  "000000100010011111",  "000000100010011011",  "000000100010010111",  "000000100010010011",  "000000100010001111",  "000000100010001011",  "000000100010000111",  "000000100010000011",  "000000100001111110",  "000000100001111010",  "000000100001110110",  "000000100001110010",  "000000100001101110",  "000000100001101001",  "000000100001100101",  "000000100001100001",  "000000100001011100",  "000000100001011000",  "000000100001010100",  "000000100001001111",  "000000100001001011",  "000000100001000110",  "000000100001000010",  "000000100000111110",  "000000100000111001",  "000000100000110101",  "000000100000110000",  "000000100000101011",  "000000100000100111",  "000000100000100010",  "000000100000011110",  "000000100000011001",  "000000100000010101",  "000000100000010000",  "000000100000001011",  "000000100000000111",  "000000100000000010",  "000000011111111101",  "000000011111111000",  "000000011111110100",  "000000011111101111",  "000000011111101010",  "000000011111100101",  "000000011111100001",  "000000011111011100",  "000000011111010111",  "000000011111010010",  "000000011111001101",  "000000011111001000",  "000000011111000011",  "000000011110111110",  "000000011110111001",  "000000011110110100",  "000000011110101111",  "000000011110101010",  "000000011110100101",  "000000011110100000",  "000000011110011011",  "000000011110010110",  "000000011110010001",  "000000011110001100",  "000000011110000111",  "000000011110000010",  "000000011101111101",  "000000011101110111",  "000000011101110010",  "000000011101101101",  "000000011101101000",  "000000011101100011",  "000000011101011101",  "000000011101011000",  "000000011101010011",  "000000011101001101",  "000000011101001000",  "000000011101000011",  "000000011100111101",  "000000011100111000",  "000000011100110011",  "000000011100101101",  "000000011100101000",  "000000011100100011",  "000000011100011101",  "000000011100011000",  "000000011100010010",  "000000011100001101",  "000000011100000111",  "000000011100000010",  "000000011011111100",  "000000011011110111",  "000000011011110001",  "000000011011101011",  "000000011011100110",  "000000011011100000",  "000000011011011011",  "000000011011010101",  "000000011011001111",  "000000011011001010",  "000000011011000100",  "000000011010111110",  "000000011010111001",  "000000011010110011",  "000000011010101101",  "000000011010100111",  "000000011010100010",  "000000011010011100",  "000000011010010110",  "000000011010010000",  "000000011010001010",  "000000011010000101",  "000000011001111111",  "000000011001111001",  "000000011001110011",  "000000011001101101",  "000000011001100111",  "000000011001100001",  "000000011001011011",  "000000011001010101",  "000000011001010000",  "000000011001001010",  "000000011001000100",  "000000011000111110",  "000000011000111000",  "000000011000110010",  "000000011000101100",  "000000011000100101",  "000000011000011111",  "000000011000011001",  "000000011000010011",  "000000011000001101",  "000000011000000111",  "000000011000000001",  "000000010111111011",  "000000010111110101",  "000000010111101111",  "000000010111101000",  "000000010111100010",  "000000010111011100",  "000000010111010110",  "000000010111010000",  "000000010111001001",  "000000010111000011",  "000000010110111101",  "000000010110110111",  "000000010110110000",  "000000010110101010",  "000000010110100100",  "000000010110011101",  "000000010110010111",  "000000010110010001",  "000000010110001010",  "000000010110000100",  "000000010101111110",  "000000010101110111",  "000000010101110001",  "000000010101101011",  "000000010101100100",  "000000010101011110",  "000000010101010111",  "000000010101010001",  "000000010101001010",  "000000010101000100",  "000000010100111101",  "000000010100110111",  "000000010100110000",  "000000010100101010",  "000000010100100011",  "000000010100011101",  "000000010100010110",  "000000010100010000",  "000000010100001001",  "000000010100000011",  "000000010011111100",  "000000010011110110",  "000000010011101111",  "000000010011101000",  "000000010011100010",  "000000010011011011",  "000000010011010101",  "000000010011001110",  "000000010011000111",  "000000010011000001",  "000000010010111010",  "000000010010110011",  "000000010010101101",  "000000010010100110",  "000000010010011111",  "000000010010011000",  "000000010010010010",  "000000010010001011",  "000000010010000100",  "000000010001111101",  "000000010001110111",  "000000010001110000",  "000000010001101001",  "000000010001100010",  "000000010001011100",  "000000010001010101",  "000000010001001110",  "000000010001000111",  "000000010001000000",  "000000010000111010",  "000000010000110011",  "000000010000101100",  "000000010000100101",  "000000010000011110",  "000000010000010111",  "000000010000010000",  "000000010000001010",  "000000010000000011",  "000000001111111100",  "000000001111110101",  "000000001111101110",  "000000001111100111",  "000000001111100000",  "000000001111011001",  "000000001111010010",  "000000001111001011",  "000000001111000100",  "000000001110111101",  "000000001110110110",  "000000001110101111",  "000000001110101000",  "000000001110100001",  "000000001110011010",  "000000001110010011",  "000000001110001100",  "000000001110000101",  "000000001101111110",  "000000001101110111",  "000000001101110000",  "000000001101101001",  "000000001101100010",  "000000001101011011",  "000000001101010100",  "000000001101001101",  "000000001101000110",  "000000001100111111",  "000000001100111000",  "000000001100110001",  "000000001100101010",  "000000001100100011",  "000000001100011100",  "000000001100010101",  "000000001100001101",  "000000001100000110",  "000000001011111111",  "000000001011111000",  "000000001011110001",  "000000001011101010",  "000000001011100011",  "000000001011011100",  "000000001011010100",  "000000001011001101",  "000000001011000110",  "000000001010111111",  "000000001010111000",  "000000001010110001",  "000000001010101001",  "000000001010100010",  "000000001010011011",  "000000001010010100",  "000000001010001101",  "000000001010000110",  "000000001001111110",  "000000001001110111",  "000000001001110000",  "000000001001101001",  "000000001001100010",  "000000001001011010",  "000000001001010011",  "000000001001001100",  "000000001001000101",  "000000001000111110",  "000000001000110110",  "000000001000101111",  "000000001000101000",  "000000001000100001",  "000000001000011001",  "000000001000010010",  "000000001000001011",  "000000001000000100",  "000000000111111100",  "000000000111110101",  "000000000111101110",  "000000000111100111",  "000000000111100000",  "000000000111011000",  "000000000111010001",  "000000000111001010",  "000000000111000010",  "000000000110111011",  "000000000110110100",  "000000000110101101",  "000000000110100101",  "000000000110011110",  "000000000110010111",  "000000000110010000",  "000000000110001000",  "000000000110000001",  "000000000101111010",  "000000000101110011",  "000000000101101011",  "000000000101100100",  "000000000101011101",  "000000000101010101",  "000000000101001110",  "000000000101000111",  "000000000101000000",  "000000000100111000",  "000000000100110001",  "000000000100101010",  "000000000100100011",  "000000000100011011",  "000000000100010100",  "000000000100001101",  "000000000100000101",  "000000000011111110",  "000000000011110111",  "000000000011110000",  "000000000011101000",  "000000000011100001",  "000000000011011010",  "000000000011010010",  "000000000011001011",  "000000000011000100",  "000000000010111101",  "000000000010110101",  "000000000010101110",  "000000000010100111",  "000000000010100000",  "000000000010011000",  "000000000010010001",  "000000000010001010",  "000000000010000010",  "000000000001111011",  "000000000001110100",  "000000000001101101",  "000000000001100101",  "000000000001011110",  "000000000001010111",  "000000000001010000",  "000000000001001000",  "000000000001000001",  "000000000000111010",  "000000000000110011",  "000000000000101011",  "000000000000100100",  "000000000000011101",  "000000000000010110",  "000000000000001110",  "000000000000000111"),("000000000000000000",  "111111111111111001",  "111111111111110010",  "111111111111101010",  "111111111111100011",  "111111111111011100",  "111111111111010101",  "111111111111001101",  "111111111111000110",  "111111111110111111",  "111111111110111000",  "111111111110110001",  "111111111110101001",  "111111111110100010",  "111111111110011011",  "111111111110010100",  "111111111110001101",  "111111111110000110",  "111111111101111110",  "111111111101110111",  "111111111101110000",  "111111111101101001",  "111111111101100010",  "111111111101011011",  "111111111101010011",  "111111111101001100",  "111111111101000101",  "111111111100111110",  "111111111100110111",  "111111111100110000",  "111111111100101001",  "111111111100100001",  "111111111100011010",  "111111111100010011",  "111111111100001100",  "111111111100000101",  "111111111011111110",  "111111111011110111",  "111111111011110000",  "111111111011101001",  "111111111011100010",  "111111111011011010",  "111111111011010011",  "111111111011001100",  "111111111011000101",  "111111111010111110",  "111111111010110111",  "111111111010110000",  "111111111010101001",  "111111111010100010",  "111111111010011011",  "111111111010010100",  "111111111010001101",  "111111111010000110",  "111111111001111111",  "111111111001111000",  "111111111001110001",  "111111111001101010",  "111111111001100011",  "111111111001011100",  "111111111001010101",  "111111111001001110",  "111111111001000111",  "111111111001000000",  "111111111000111001",  "111111111000110010",  "111111111000101100",  "111111111000100101",  "111111111000011110",  "111111111000010111",  "111111111000010000",  "111111111000001001",  "111111111000000010",  "111111110111111011",  "111111110111110100",  "111111110111101110",  "111111110111100111",  "111111110111100000",  "111111110111011001",  "111111110111010010",  "111111110111001011",  "111111110111000101",  "111111110110111110",  "111111110110110111",  "111111110110110000",  "111111110110101001",  "111111110110100011",  "111111110110011100",  "111111110110010101",  "111111110110001110",  "111111110110001000",  "111111110110000001",  "111111110101111010",  "111111110101110011",  "111111110101101101",  "111111110101100110",  "111111110101011111",  "111111110101011001",  "111111110101010010",  "111111110101001011",  "111111110101000101",  "111111110100111110",  "111111110100110111",  "111111110100110001",  "111111110100101010",  "111111110100100100",  "111111110100011101",  "111111110100010110",  "111111110100010000",  "111111110100001001",  "111111110100000011",  "111111110011111100",  "111111110011110110",  "111111110011101111",  "111111110011101000",  "111111110011100010",  "111111110011011011",  "111111110011010101",  "111111110011001110",  "111111110011001000",  "111111110011000010",  "111111110010111011",  "111111110010110101",  "111111110010101110",  "111111110010101000",  "111111110010100001",  "111111110010011011",  "111111110010010101",  "111111110010001110",  "111111110010001000",  "111111110010000001",  "111111110001111011",  "111111110001110101",  "111111110001101110",  "111111110001101000",  "111111110001100010",  "111111110001011100",  "111111110001010101",  "111111110001001111",  "111111110001001001",  "111111110001000010",  "111111110000111100",  "111111110000110110",  "111111110000110000",  "111111110000101010",  "111111110000100011",  "111111110000011101",  "111111110000010111",  "111111110000010001",  "111111110000001011",  "111111110000000101",  "111111101111111110",  "111111101111111000",  "111111101111110010",  "111111101111101100",  "111111101111100110",  "111111101111100000",  "111111101111011010",  "111111101111010100",  "111111101111001110",  "111111101111001000",  "111111101111000010",  "111111101110111100",  "111111101110110110",  "111111101110110000",  "111111101110101010",  "111111101110100100",  "111111101110011110",  "111111101110011000",  "111111101110010010",  "111111101110001100",  "111111101110000111",  "111111101110000001",  "111111101101111011",  "111111101101110101",  "111111101101101111",  "111111101101101001",  "111111101101100100",  "111111101101011110",  "111111101101011000",  "111111101101010010",  "111111101101001100",  "111111101101000111",  "111111101101000001",  "111111101100111011",  "111111101100110110",  "111111101100110000",  "111111101100101010",  "111111101100100101",  "111111101100011111",  "111111101100011001",  "111111101100010100",  "111111101100001110",  "111111101100001001",  "111111101100000011",  "111111101011111101",  "111111101011111000",  "111111101011110010",  "111111101011101101",  "111111101011100111",  "111111101011100010",  "111111101011011100",  "111111101011010111",  "111111101011010010",  "111111101011001100",  "111111101011000111",  "111111101011000001",  "111111101010111100",  "111111101010110111",  "111111101010110001",  "111111101010101100",  "111111101010100111",  "111111101010100001",  "111111101010011100",  "111111101010010111",  "111111101010010001",  "111111101010001100",  "111111101010000111",  "111111101010000010",  "111111101001111100",  "111111101001110111",  "111111101001110010",  "111111101001101101",  "111111101001101000",  "111111101001100011",  "111111101001011110",  "111111101001011000",  "111111101001010011",  "111111101001001110",  "111111101001001001",  "111111101001000100",  "111111101000111111",  "111111101000111010",  "111111101000110101",  "111111101000110000",  "111111101000101011",  "111111101000100110",  "111111101000100001",  "111111101000011101",  "111111101000011000",  "111111101000010011",  "111111101000001110",  "111111101000001001",  "111111101000000100",  "111111100111111111",  "111111100111111011",  "111111100111110110",  "111111100111110001",  "111111100111101100",  "111111100111101000",  "111111100111100011",  "111111100111011110",  "111111100111011010",  "111111100111010101",  "111111100111010000",  "111111100111001100",  "111111100111000111",  "111111100111000010",  "111111100110111110",  "111111100110111001",  "111111100110110101",  "111111100110110000",  "111111100110101100",  "111111100110100111",  "111111100110100011",  "111111100110011110",  "111111100110011010",  "111111100110010101",  "111111100110010001",  "111111100110001101",  "111111100110001000",  "111111100110000100",  "111111100101111111",  "111111100101111011",  "111111100101110111",  "111111100101110011",  "111111100101101110",  "111111100101101010",  "111111100101100110",  "111111100101100010",  "111111100101011101",  "111111100101011001",  "111111100101010101",  "111111100101010001",  "111111100101001101",  "111111100101001001",  "111111100101000100",  "111111100101000000",  "111111100100111100",  "111111100100111000",  "111111100100110100",  "111111100100110000",  "111111100100101100",  "111111100100101000",  "111111100100100100",  "111111100100100000",  "111111100100011100",  "111111100100011001",  "111111100100010101",  "111111100100010001",  "111111100100001101",  "111111100100001001",  "111111100100000101",  "111111100100000001",  "111111100011111110",  "111111100011111010",  "111111100011110110",  "111111100011110011",  "111111100011101111",  "111111100011101011",  "111111100011100111",  "111111100011100100",  "111111100011100000",  "111111100011011101",  "111111100011011001",  "111111100011010101",  "111111100011010010",  "111111100011001110",  "111111100011001011",  "111111100011000111",  "111111100011000100",  "111111100011000000",  "111111100010111101",  "111111100010111001",  "111111100010110110",  "111111100010110011",  "111111100010101111",  "111111100010101100",  "111111100010101001",  "111111100010100101",  "111111100010100010",  "111111100010011111",  "111111100010011100",  "111111100010011000",  "111111100010010101",  "111111100010010010",  "111111100010001111",  "111111100010001100",  "111111100010001000",  "111111100010000101",  "111111100010000010",  "111111100001111111",  "111111100001111100",  "111111100001111001",  "111111100001110110",  "111111100001110011",  "111111100001110000",  "111111100001101101",  "111111100001101010",  "111111100001100111",  "111111100001100100",  "111111100001100001",  "111111100001011110",  "111111100001011100",  "111111100001011001",  "111111100001010110",  "111111100001010011",  "111111100001010000",  "111111100001001110",  "111111100001001011",  "111111100001001000",  "111111100001000110",  "111111100001000011",  "111111100001000000",  "111111100000111110",  "111111100000111011",  "111111100000111000",  "111111100000110110",  "111111100000110011",  "111111100000110001",  "111111100000101110",  "111111100000101100",  "111111100000101001",  "111111100000100111",  "111111100000100100",  "111111100000100010",  "111111100000100000",  "111111100000011101",  "111111100000011011",  "111111100000011000",  "111111100000010110",  "111111100000010100",  "111111100000010010",  "111111100000001111",  "111111100000001101",  "111111100000001011",  "111111100000001001",  "111111100000000110",  "111111100000000100",  "111111100000000010",  "111111100000000000",  "111111011111111110",  "111111011111111100",  "111111011111111010",  "111111011111111000",  "111111011111110110",  "111111011111110100",  "111111011111110010",  "111111011111110000",  "111111011111101110",  "111111011111101100",  "111111011111101010",  "111111011111101000",  "111111011111100110",  "111111011111100101",  "111111011111100011",  "111111011111100001",  "111111011111011111",  "111111011111011101",  "111111011111011100",  "111111011111011010",  "111111011111011000",  "111111011111010111",  "111111011111010101",  "111111011111010011",  "111111011111010010",  "111111011111010000",  "111111011111001111",  "111111011111001101",  "111111011111001011",  "111111011111001010",  "111111011111001000",  "111111011111000111",  "111111011111000110",  "111111011111000100",  "111111011111000011",  "111111011111000001",  "111111011111000000",  "111111011110111111",  "111111011110111101",  "111111011110111100",  "111111011110111011",  "111111011110111001",  "111111011110111000",  "111111011110110111",  "111111011110110110",  "111111011110110101",  "111111011110110011",  "111111011110110010",  "111111011110110001",  "111111011110110000",  "111111011110101111",  "111111011110101110",  "111111011110101101",  "111111011110101100",  "111111011110101011",  "111111011110101010",  "111111011110101001",  "111111011110101000",  "111111011110100111",  "111111011110100110",  "111111011110100101",  "111111011110100100",  "111111011110100100",  "111111011110100011",  "111111011110100010",  "111111011110100001",  "111111011110100001",  "111111011110100000",  "111111011110011111",  "111111011110011110",  "111111011110011110",  "111111011110011101",  "111111011110011100",  "111111011110011100",  "111111011110011011",  "111111011110011011",  "111111011110011010",  "111111011110011010",  "111111011110011001",  "111111011110011001",  "111111011110011000",  "111111011110011000",  "111111011110010111",  "111111011110010111",  "111111011110010110",  "111111011110010110",  "111111011110010110",  "111111011110010101",  "111111011110010101",  "111111011110010101",  "111111011110010101",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010011",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010100",  "111111011110010101",  "111111011110010101",  "111111011110010101",  "111111011110010110",  "111111011110010110",  "111111011110010110",  "111111011110010111",  "111111011110010111",  "111111011110010111",  "111111011110011000",  "111111011110011000",  "111111011110011001",  "111111011110011001",  "111111011110011010",  "111111011110011010",  "111111011110011011",  "111111011110011011",  "111111011110011100",  "111111011110011101",  "111111011110011101",  "111111011110011110",  "111111011110011111",  "111111011110011111",  "111111011110100000",  "111111011110100001",  "111111011110100010",  "111111011110100010",  "111111011110100011",  "111111011110100100",  "111111011110100101",  "111111011110100110",  "111111011110100110",  "111111011110100111",  "111111011110101000",  "111111011110101001",  "111111011110101010",  "111111011110101011",  "111111011110101100",  "111111011110101101",  "111111011110101110",  "111111011110101111",  "111111011110110000",  "111111011110110001",  "111111011110110010",  "111111011110110100",  "111111011110110101",  "111111011110110110",  "111111011110110111",  "111111011110111000",  "111111011110111010",  "111111011110111011",  "111111011110111100",  "111111011110111101",  "111111011110111111",  "111111011111000000",  "111111011111000001",  "111111011111000011",  "111111011111000100",  "111111011111000101",  "111111011111000111",  "111111011111001000",  "111111011111001010",  "111111011111001011",  "111111011111001101",  "111111011111001110",  "111111011111010000",  "111111011111010001",  "111111011111010011",  "111111011111010101",  "111111011111010110",  "111111011111011000",  "111111011111011001",  "111111011111011011",  "111111011111011101",  "111111011111011111",  "111111011111100000",  "111111011111100010",  "111111011111100100",  "111111011111100110",  "111111011111100111",  "111111011111101001",  "111111011111101011",  "111111011111101101",  "111111011111101111",  "111111011111110001",  "111111011111110011",  "111111011111110101",  "111111011111110110",  "111111011111111000",  "111111011111111010",  "111111011111111100",  "111111011111111110",  "111111100000000001",  "111111100000000011",  "111111100000000101",  "111111100000000111",  "111111100000001001",  "111111100000001011",  "111111100000001101",  "111111100000001111",  "111111100000010010",  "111111100000010100",  "111111100000010110",  "111111100000011000",  "111111100000011011",  "111111100000011101",  "111111100000011111",  "111111100000100010",  "111111100000100100",  "111111100000100110",  "111111100000101001",  "111111100000101011",  "111111100000101101",  "111111100000110000",  "111111100000110010",  "111111100000110101",  "111111100000110111",  "111111100000111010",  "111111100000111100",  "111111100000111111",  "111111100001000001",  "111111100001000100",  "111111100001000111",  "111111100001001001",  "111111100001001100",  "111111100001001110",  "111111100001010001",  "111111100001010100",  "111111100001010111",  "111111100001011001",  "111111100001011100",  "111111100001011111",  "111111100001100001",  "111111100001100100",  "111111100001100111",  "111111100001101010",  "111111100001101101",  "111111100001110000",  "111111100001110010",  "111111100001110101",  "111111100001111000",  "111111100001111011",  "111111100001111110",  "111111100010000001",  "111111100010000100",  "111111100010000111",  "111111100010001010",  "111111100010001101",  "111111100010010000",  "111111100010010011",  "111111100010010110",  "111111100010011001",  "111111100010011101",  "111111100010100000",  "111111100010100011",  "111111100010100110",  "111111100010101001",  "111111100010101100",  "111111100010110000",  "111111100010110011",  "111111100010110110",  "111111100010111001",  "111111100010111101",  "111111100011000000",  "111111100011000011",  "111111100011000111",  "111111100011001010",  "111111100011001101",  "111111100011010001",  "111111100011010100",  "111111100011010111",  "111111100011011011",  "111111100011011110",  "111111100011100010",  "111111100011100101",  "111111100011101001",  "111111100011101100",  "111111100011110000",  "111111100011110011",  "111111100011110111",  "111111100011111010",  "111111100011111110",  "111111100100000010",  "111111100100000101",  "111111100100001001",  "111111100100001101",  "111111100100010000",  "111111100100010100",  "111111100100011000",  "111111100100011011",  "111111100100011111",  "111111100100100011",  "111111100100100110",  "111111100100101010",  "111111100100101110",  "111111100100110010",  "111111100100110110",  "111111100100111001",  "111111100100111101",  "111111100101000001",  "111111100101000101",  "111111100101001001",  "111111100101001101",  "111111100101010001",  "111111100101010101",  "111111100101011001",  "111111100101011101",  "111111100101100001",  "111111100101100101",  "111111100101101001",  "111111100101101101",  "111111100101110001",  "111111100101110101",  "111111100101111001",  "111111100101111101",  "111111100110000001",  "111111100110000101",  "111111100110001001",  "111111100110001101",  "111111100110010010",  "111111100110010110",  "111111100110011010",  "111111100110011110",  "111111100110100010",  "111111100110100110",  "111111100110101011",  "111111100110101111",  "111111100110110011",  "111111100110111000",  "111111100110111100",  "111111100111000000",  "111111100111000100",  "111111100111001001",  "111111100111001101",  "111111100111010001",  "111111100111010110",  "111111100111011010",  "111111100111011111",  "111111100111100011",  "111111100111100111",  "111111100111101100",  "111111100111110000",  "111111100111110101",  "111111100111111001",  "111111100111111110",  "111111101000000010",  "111111101000000111",  "111111101000001011",  "111111101000010000",  "111111101000010100",  "111111101000011001",  "111111101000011110",  "111111101000100010",  "111111101000100111",  "111111101000101011",  "111111101000110000",  "111111101000110101",  "111111101000111001",  "111111101000111110",  "111111101001000011",  "111111101001000111",  "111111101001001100",  "111111101001010001",  "111111101001010110",  "111111101001011010",  "111111101001011111",  "111111101001100100",  "111111101001101001",  "111111101001101101",  "111111101001110010",  "111111101001110111",  "111111101001111100",  "111111101010000001",  "111111101010000101",  "111111101010001010",  "111111101010001111",  "111111101010010100",  "111111101010011001",  "111111101010011110",  "111111101010100011",  "111111101010101000",  "111111101010101101",  "111111101010110010",  "111111101010110111",  "111111101010111100",  "111111101011000000",  "111111101011000101",  "111111101011001010",  "111111101011010000",  "111111101011010101",  "111111101011011010",  "111111101011011111",  "111111101011100100",  "111111101011101001",  "111111101011101110",  "111111101011110011",  "111111101011111000",  "111111101011111101",  "111111101100000010",  "111111101100000111",  "111111101100001100",  "111111101100010010",  "111111101100010111",  "111111101100011100",  "111111101100100001",  "111111101100100110",  "111111101100101100",  "111111101100110001",  "111111101100110110",  "111111101100111011",  "111111101101000000",  "111111101101000110",  "111111101101001011",  "111111101101010000",  "111111101101010101",  "111111101101011011",  "111111101101100000",  "111111101101100101",  "111111101101101011",  "111111101101110000",  "111111101101110101",  "111111101101111011",  "111111101110000000",  "111111101110000101",  "111111101110001011",  "111111101110010000",  "111111101110010110",  "111111101110011011",  "111111101110100000",  "111111101110100110",  "111111101110101011",  "111111101110110001",  "111111101110110110",  "111111101110111011",  "111111101111000001",  "111111101111000110",  "111111101111001100",  "111111101111010001",  "111111101111010111",  "111111101111011100",  "111111101111100010",  "111111101111100111",  "111111101111101101",  "111111101111110010",  "111111101111111000",  "111111101111111101",  "111111110000000011",  "111111110000001001",  "111111110000001110",  "111111110000010100",  "111111110000011001",  "111111110000011111",  "111111110000100101",  "111111110000101010",  "111111110000110000",  "111111110000110101",  "111111110000111011",  "111111110001000001",  "111111110001000110",  "111111110001001100",  "111111110001010010",  "111111110001010111",  "111111110001011101",  "111111110001100011",  "111111110001101000",  "111111110001101110",  "111111110001110100",  "111111110001111001",  "111111110001111111",  "111111110010000101",  "111111110010001010",  "111111110010010000",  "111111110010010110",  "111111110010011100",  "111111110010100001",  "111111110010100111",  "111111110010101101",  "111111110010110011",  "111111110010111000",  "111111110010111110",  "111111110011000100",  "111111110011001010",  "111111110011010000",  "111111110011010101",  "111111110011011011",  "111111110011100001",  "111111110011100111",  "111111110011101101",  "111111110011110010",  "111111110011111000",  "111111110011111110",  "111111110100000100",  "111111110100001010",  "111111110100010000",  "111111110100010110",  "111111110100011011",  "111111110100100001",  "111111110100100111",  "111111110100101101",  "111111110100110011",  "111111110100111001",  "111111110100111111",  "111111110101000101",  "111111110101001010",  "111111110101010000",  "111111110101010110",  "111111110101011100",  "111111110101100010",  "111111110101101000",  "111111110101101110",  "111111110101110100",  "111111110101111010",  "111111110110000000",  "111111110110000110",  "111111110110001100",  "111111110110010010",  "111111110110011000",  "111111110110011101",  "111111110110100011",  "111111110110101001",  "111111110110101111",  "111111110110110101",  "111111110110111011",  "111111110111000001",  "111111110111000111",  "111111110111001101",  "111111110111010011",  "111111110111011001",  "111111110111011111",  "111111110111100101",  "111111110111101011",  "111111110111110001",  "111111110111110111",  "111111110111111101",  "111111111000000011",  "111111111000001001",  "111111111000001111",  "111111111000010101",  "111111111000011011",  "111111111000100001",  "111111111000100111",  "111111111000101101",  "111111111000110011",  "111111111000111001",  "111111111000111111",  "111111111001000110",  "111111111001001100",  "111111111001010010",  "111111111001011000",  "111111111001011110",  "111111111001100100",  "111111111001101010",  "111111111001110000",  "111111111001110110",  "111111111001111100",  "111111111010000010",  "111111111010001000",  "111111111010001110",  "111111111010010100",  "111111111010011010",  "111111111010100000",  "111111111010100110",  "111111111010101100",  "111111111010110010",  "111111111010111001",  "111111111010111111",  "111111111011000101",  "111111111011001011",  "111111111011010001",  "111111111011010111",  "111111111011011101",  "111111111011100011",  "111111111011101001",  "111111111011101111",  "111111111011110101",  "111111111011111011",  "111111111100000001",  "111111111100000111",  "111111111100001110",  "111111111100010100",  "111111111100011010",  "111111111100100000",  "111111111100100110",  "111111111100101100",  "111111111100110010",  "111111111100111000",  "111111111100111110",  "111111111101000100",  "111111111101001010",  "111111111101010000",  "111111111101010110",  "111111111101011101",  "111111111101100011",  "111111111101101001",  "111111111101101111",  "111111111101110101",  "111111111101111011",  "111111111110000001",  "111111111110000111",  "111111111110001101",  "111111111110010011",  "111111111110011001",  "111111111110011111",  "111111111110100101",  "111111111110101011",  "111111111110110001",  "111111111110110111",  "111111111110111110",  "111111111111000100",  "111111111111001010",  "111111111111010000",  "111111111111010110",  "111111111111011100",  "111111111111100010",  "111111111111101000",  "111111111111101110",  "111111111111110100",  "111111111111111010"),("000000000000000000",  "000000000000000110",  "000000000000001100",  "000000000000010010",  "000000000000011000",  "000000000000011110",  "000000000000100100",  "000000000000101010",  "000000000000110000",  "000000000000110110",  "000000000000111100",  "000000000001000010",  "000000000001001000",  "000000000001001110",  "000000000001010100",  "000000000001011010",  "000000000001100000",  "000000000001100110",  "000000000001101100",  "000000000001110010",  "000000000001111000",  "000000000001111110",  "000000000010000100",  "000000000010001010",  "000000000010010000",  "000000000010010110",  "000000000010011100",  "000000000010100010",  "000000000010101000",  "000000000010101110",  "000000000010110100",  "000000000010111010",  "000000000011000000",  "000000000011000110",  "000000000011001100",  "000000000011010001",  "000000000011010111",  "000000000011011101",  "000000000011100011",  "000000000011101001",  "000000000011101111",  "000000000011110101",  "000000000011111011",  "000000000100000001",  "000000000100000111",  "000000000100001100",  "000000000100010010",  "000000000100011000",  "000000000100011110",  "000000000100100100",  "000000000100101010",  "000000000100110000",  "000000000100110110",  "000000000100111011",  "000000000101000001",  "000000000101000111",  "000000000101001101",  "000000000101010011",  "000000000101011001",  "000000000101011110",  "000000000101100100",  "000000000101101010",  "000000000101110000",  "000000000101110110",  "000000000101111011",  "000000000110000001",  "000000000110000111",  "000000000110001101",  "000000000110010010",  "000000000110011000",  "000000000110011110",  "000000000110100100",  "000000000110101001",  "000000000110101111",  "000000000110110101",  "000000000110111011",  "000000000111000000",  "000000000111000110",  "000000000111001100",  "000000000111010001",  "000000000111010111",  "000000000111011101",  "000000000111100010",  "000000000111101000",  "000000000111101110",  "000000000111110011",  "000000000111111001",  "000000000111111111",  "000000001000000100",  "000000001000001010",  "000000001000010000",  "000000001000010101",  "000000001000011011",  "000000001000100000",  "000000001000100110",  "000000001000101100",  "000000001000110001",  "000000001000110111",  "000000001000111100",  "000000001001000010",  "000000001001000111",  "000000001001001101",  "000000001001010011",  "000000001001011000",  "000000001001011110",  "000000001001100011",  "000000001001101001",  "000000001001101110",  "000000001001110100",  "000000001001111001",  "000000001001111111",  "000000001010000100",  "000000001010001001",  "000000001010001111",  "000000001010010100",  "000000001010011010",  "000000001010011111",  "000000001010100101",  "000000001010101010",  "000000001010101111",  "000000001010110101",  "000000001010111010",  "000000001011000000",  "000000001011000101",  "000000001011001010",  "000000001011010000",  "000000001011010101",  "000000001011011010",  "000000001011100000",  "000000001011100101",  "000000001011101010",  "000000001011110000",  "000000001011110101",  "000000001011111010",  "000000001011111111",  "000000001100000101",  "000000001100001010",  "000000001100001111",  "000000001100010100",  "000000001100011010",  "000000001100011111",  "000000001100100100",  "000000001100101001",  "000000001100101110",  "000000001100110100",  "000000001100111001",  "000000001100111110",  "000000001101000011",  "000000001101001000",  "000000001101001101",  "000000001101010010",  "000000001101011000",  "000000001101011101",  "000000001101100010",  "000000001101100111",  "000000001101101100",  "000000001101110001",  "000000001101110110",  "000000001101111011",  "000000001110000000",  "000000001110000101",  "000000001110001010",  "000000001110001111",  "000000001110010100",  "000000001110011001",  "000000001110011110",  "000000001110100011",  "000000001110101000",  "000000001110101101",  "000000001110110010",  "000000001110110111",  "000000001110111100",  "000000001111000000",  "000000001111000101",  "000000001111001010",  "000000001111001111",  "000000001111010100",  "000000001111011001",  "000000001111011110",  "000000001111100010",  "000000001111100111",  "000000001111101100",  "000000001111110001",  "000000001111110101",  "000000001111111010",  "000000001111111111",  "000000010000000100",  "000000010000001000",  "000000010000001101",  "000000010000010010",  "000000010000010111",  "000000010000011011",  "000000010000100000",  "000000010000100101",  "000000010000101001",  "000000010000101110",  "000000010000110010",  "000000010000110111",  "000000010000111100",  "000000010001000000",  "000000010001000101",  "000000010001001001",  "000000010001001110",  "000000010001010010",  "000000010001010111",  "000000010001011011",  "000000010001100000",  "000000010001100100",  "000000010001101001",  "000000010001101101",  "000000010001110010",  "000000010001110110",  "000000010001111011",  "000000010001111111",  "000000010010000100",  "000000010010001000",  "000000010010001100",  "000000010010010001",  "000000010010010101",  "000000010010011001",  "000000010010011110",  "000000010010100010",  "000000010010100110",  "000000010010101011",  "000000010010101111",  "000000010010110011",  "000000010010110111",  "000000010010111100",  "000000010011000000",  "000000010011000100",  "000000010011001000",  "000000010011001100",  "000000010011010001",  "000000010011010101",  "000000010011011001",  "000000010011011101",  "000000010011100001",  "000000010011100101",  "000000010011101001",  "000000010011101101",  "000000010011110001",  "000000010011110101",  "000000010011111010",  "000000010011111110",  "000000010100000010",  "000000010100000110",  "000000010100001010",  "000000010100001110",  "000000010100010001",  "000000010100010101",  "000000010100011001",  "000000010100011101",  "000000010100100001",  "000000010100100101",  "000000010100101001",  "000000010100101101",  "000000010100110001",  "000000010100110100",  "000000010100111000",  "000000010100111100",  "000000010101000000",  "000000010101000100",  "000000010101000111",  "000000010101001011",  "000000010101001111",  "000000010101010011",  "000000010101010110",  "000000010101011010",  "000000010101011110",  "000000010101100001",  "000000010101100101",  "000000010101101001",  "000000010101101100",  "000000010101110000",  "000000010101110011",  "000000010101110111",  "000000010101111011",  "000000010101111110",  "000000010110000010",  "000000010110000101",  "000000010110001001",  "000000010110001100",  "000000010110010000",  "000000010110010011",  "000000010110010111",  "000000010110011010",  "000000010110011101",  "000000010110100001",  "000000010110100100",  "000000010110101000",  "000000010110101011",  "000000010110101110",  "000000010110110010",  "000000010110110101",  "000000010110111000",  "000000010110111011",  "000000010110111111",  "000000010111000010",  "000000010111000101",  "000000010111001000",  "000000010111001100",  "000000010111001111",  "000000010111010010",  "000000010111010101",  "000000010111011000",  "000000010111011011",  "000000010111011111",  "000000010111100010",  "000000010111100101",  "000000010111101000",  "000000010111101011",  "000000010111101110",  "000000010111110001",  "000000010111110100",  "000000010111110111",  "000000010111111010",  "000000010111111101",  "000000011000000000",  "000000011000000011",  "000000011000000110",  "000000011000001001",  "000000011000001011",  "000000011000001110",  "000000011000010001",  "000000011000010100",  "000000011000010111",  "000000011000011010",  "000000011000011100",  "000000011000011111",  "000000011000100010",  "000000011000100101",  "000000011000100111",  "000000011000101010",  "000000011000101101",  "000000011000101111",  "000000011000110010",  "000000011000110101",  "000000011000110111",  "000000011000111010",  "000000011000111101",  "000000011000111111",  "000000011001000010",  "000000011001000100",  "000000011001000111",  "000000011001001001",  "000000011001001100",  "000000011001001110",  "000000011001010001",  "000000011001010011",  "000000011001010110",  "000000011001011000",  "000000011001011011",  "000000011001011101",  "000000011001011111",  "000000011001100010",  "000000011001100100",  "000000011001100110",  "000000011001101001",  "000000011001101011",  "000000011001101101",  "000000011001101111",  "000000011001110010",  "000000011001110100",  "000000011001110110",  "000000011001111000",  "000000011001111010",  "000000011001111101",  "000000011001111111",  "000000011010000001",  "000000011010000011",  "000000011010000101",  "000000011010000111",  "000000011010001001",  "000000011010001011",  "000000011010001101",  "000000011010001111",  "000000011010010001",  "000000011010010011",  "000000011010010101",  "000000011010010111",  "000000011010011001",  "000000011010011011",  "000000011010011101",  "000000011010011111",  "000000011010100001",  "000000011010100011",  "000000011010100100",  "000000011010100110",  "000000011010101000",  "000000011010101010",  "000000011010101100",  "000000011010101101",  "000000011010101111",  "000000011010110001",  "000000011010110010",  "000000011010110100",  "000000011010110110",  "000000011010110111",  "000000011010111001",  "000000011010111011",  "000000011010111100",  "000000011010111110",  "000000011010111111",  "000000011011000001",  "000000011011000010",  "000000011011000100",  "000000011011000101",  "000000011011000111",  "000000011011001000",  "000000011011001010",  "000000011011001011",  "000000011011001101",  "000000011011001110",  "000000011011001111",  "000000011011010001",  "000000011011010010",  "000000011011010011",  "000000011011010101",  "000000011011010110",  "000000011011010111",  "000000011011011001",  "000000011011011010",  "000000011011011011",  "000000011011011100",  "000000011011011101",  "000000011011011111",  "000000011011100000",  "000000011011100001",  "000000011011100010",  "000000011011100011",  "000000011011100100",  "000000011011100101",  "000000011011100110",  "000000011011100111",  "000000011011101000",  "000000011011101001",  "000000011011101010",  "000000011011101011",  "000000011011101100",  "000000011011101101",  "000000011011101110",  "000000011011101111",  "000000011011110000",  "000000011011110001",  "000000011011110001",  "000000011011110010",  "000000011011110011",  "000000011011110100",  "000000011011110101",  "000000011011110101",  "000000011011110110",  "000000011011110111",  "000000011011111000",  "000000011011111000",  "000000011011111001",  "000000011011111010",  "000000011011111010",  "000000011011111011",  "000000011011111100",  "000000011011111100",  "000000011011111101",  "000000011011111101",  "000000011011111110",  "000000011011111110",  "000000011011111111",  "000000011011111111",  "000000011100000000",  "000000011100000000",  "000000011100000001",  "000000011100000001",  "000000011100000001",  "000000011100000010",  "000000011100000010",  "000000011100000011",  "000000011100000011",  "000000011100000011",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000110",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000101",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000100",  "000000011100000011",  "000000011100000011",  "000000011100000011",  "000000011100000010",  "000000011100000010",  "000000011100000001",  "000000011100000001",  "000000011100000001",  "000000011100000000",  "000000011100000000",  "000000011011111111",  "000000011011111111",  "000000011011111110",  "000000011011111110",  "000000011011111101",  "000000011011111101",  "000000011011111100",  "000000011011111100",  "000000011011111011",  "000000011011111010",  "000000011011111010",  "000000011011111001",  "000000011011111000",  "000000011011111000",  "000000011011110111",  "000000011011110110",  "000000011011110110",  "000000011011110101",  "000000011011110100",  "000000011011110011",  "000000011011110011",  "000000011011110010",  "000000011011110001",  "000000011011110000",  "000000011011101111",  "000000011011101110",  "000000011011101101",  "000000011011101100",  "000000011011101100",  "000000011011101011",  "000000011011101010",  "000000011011101001",  "000000011011101000",  "000000011011100111",  "000000011011100110",  "000000011011100101",  "000000011011100100",  "000000011011100010",  "000000011011100001",  "000000011011100000",  "000000011011011111",  "000000011011011110",  "000000011011011101",  "000000011011011100",  "000000011011011010",  "000000011011011001",  "000000011011011000",  "000000011011010111",  "000000011011010110",  "000000011011010100",  "000000011011010011",  "000000011011010010",  "000000011011010000",  "000000011011001111",  "000000011011001110",  "000000011011001100",  "000000011011001011",  "000000011011001010",  "000000011011001000",  "000000011011000111",  "000000011011000101",  "000000011011000100",  "000000011011000010",  "000000011011000001",  "000000011010111111",  "000000011010111110",  "000000011010111100",  "000000011010111011",  "000000011010111001",  "000000011010111000",  "000000011010110110",  "000000011010110100",  "000000011010110011",  "000000011010110001",  "000000011010101111",  "000000011010101110",  "000000011010101100",  "000000011010101010",  "000000011010101001",  "000000011010100111",  "000000011010100101",  "000000011010100011",  "000000011010100001",  "000000011010100000",  "000000011010011110",  "000000011010011100",  "000000011010011010",  "000000011010011000",  "000000011010010110",  "000000011010010101",  "000000011010010011",  "000000011010010001",  "000000011010001111",  "000000011010001101",  "000000011010001011",  "000000011010001001",  "000000011010000111",  "000000011010000101",  "000000011010000011",  "000000011010000001",  "000000011001111111",  "000000011001111101",  "000000011001111010",  "000000011001111000",  "000000011001110110",  "000000011001110100",  "000000011001110010",  "000000011001110000",  "000000011001101110",  "000000011001101011",  "000000011001101001",  "000000011001100111",  "000000011001100101",  "000000011001100010",  "000000011001100000",  "000000011001011110",  "000000011001011100",  "000000011001011001",  "000000011001010111",  "000000011001010101",  "000000011001010010",  "000000011001010000",  "000000011001001110",  "000000011001001011",  "000000011001001001",  "000000011001000110",  "000000011001000100",  "000000011001000001",  "000000011000111111",  "000000011000111100",  "000000011000111010",  "000000011000110111",  "000000011000110101",  "000000011000110010",  "000000011000110000",  "000000011000101101",  "000000011000101011",  "000000011000101000",  "000000011000100101",  "000000011000100011",  "000000011000100000",  "000000011000011101",  "000000011000011011",  "000000011000011000",  "000000011000010101",  "000000011000010011",  "000000011000010000",  "000000011000001101",  "000000011000001011",  "000000011000001000",  "000000011000000101",  "000000011000000010",  "000000010111111111",  "000000010111111101",  "000000010111111010",  "000000010111110111",  "000000010111110100",  "000000010111110001",  "000000010111101110",  "000000010111101011",  "000000010111101000",  "000000010111100110",  "000000010111100011",  "000000010111100000",  "000000010111011101",  "000000010111011010",  "000000010111010111",  "000000010111010100",  "000000010111010001",  "000000010111001110",  "000000010111001011",  "000000010111001000",  "000000010111000100",  "000000010111000001",  "000000010110111110",  "000000010110111011",  "000000010110111000",  "000000010110110101",  "000000010110110010",  "000000010110101111",  "000000010110101011",  "000000010110101000",  "000000010110100101",  "000000010110100010",  "000000010110011111",  "000000010110011011",  "000000010110011000",  "000000010110010101",  "000000010110010010",  "000000010110001110",  "000000010110001011",  "000000010110001000",  "000000010110000100",  "000000010110000001",  "000000010101111110",  "000000010101111010",  "000000010101110111",  "000000010101110100",  "000000010101110000",  "000000010101101101",  "000000010101101001",  "000000010101100110",  "000000010101100011",  "000000010101011111",  "000000010101011100",  "000000010101011000",  "000000010101010101",  "000000010101010001",  "000000010101001110",  "000000010101001010",  "000000010101000111",  "000000010101000011",  "000000010101000000",  "000000010100111100",  "000000010100111000",  "000000010100110101",  "000000010100110001",  "000000010100101110",  "000000010100101010",  "000000010100100110",  "000000010100100011",  "000000010100011111",  "000000010100011011",  "000000010100011000",  "000000010100010100",  "000000010100010000",  "000000010100001101",  "000000010100001001",  "000000010100000101",  "000000010100000001",  "000000010011111110",  "000000010011111010",  "000000010011110110",  "000000010011110010",  "000000010011101110",  "000000010011101011",  "000000010011100111",  "000000010011100011",  "000000010011011111",  "000000010011011011",  "000000010011010111",  "000000010011010100",  "000000010011010000",  "000000010011001100",  "000000010011001000",  "000000010011000100",  "000000010011000000",  "000000010010111100",  "000000010010111000",  "000000010010110100",  "000000010010110000",  "000000010010101100",  "000000010010101000",  "000000010010100100",  "000000010010100000",  "000000010010011100",  "000000010010011000",  "000000010010010100",  "000000010010010000",  "000000010010001100",  "000000010010001000",  "000000010010000100",  "000000010010000000",  "000000010001111100",  "000000010001111000",  "000000010001110100",  "000000010001110000",  "000000010001101011",  "000000010001100111",  "000000010001100011",  "000000010001011111",  "000000010001011011",  "000000010001010111",  "000000010001010011",  "000000010001001110",  "000000010001001010",  "000000010001000110",  "000000010001000010",  "000000010000111110",  "000000010000111001",  "000000010000110101",  "000000010000110001",  "000000010000101101",  "000000010000101000",  "000000010000100100",  "000000010000100000",  "000000010000011011",  "000000010000010111",  "000000010000010011",  "000000010000001110",  "000000010000001010",  "000000010000000110",  "000000010000000001",  "000000001111111101",  "000000001111111001",  "000000001111110100",  "000000001111110000",  "000000001111101100",  "000000001111100111",  "000000001111100011",  "000000001111011110",  "000000001111011010",  "000000001111010110",  "000000001111010001",  "000000001111001101",  "000000001111001000",  "000000001111000100",  "000000001110111111",  "000000001110111011",  "000000001110110110",  "000000001110110010",  "000000001110101101",  "000000001110101001",  "000000001110100100",  "000000001110100000",  "000000001110011011",  "000000001110010111",  "000000001110010010",  "000000001110001110",  "000000001110001001",  "000000001110000101",  "000000001110000000",  "000000001101111100",  "000000001101110111",  "000000001101110010",  "000000001101101110",  "000000001101101001",  "000000001101100101",  "000000001101100000",  "000000001101011011",  "000000001101010111",  "000000001101010010",  "000000001101001110",  "000000001101001001",  "000000001101000100",  "000000001101000000",  "000000001100111011",  "000000001100110110",  "000000001100110010",  "000000001100101101",  "000000001100101000",  "000000001100100100",  "000000001100011111",  "000000001100011010",  "000000001100010110",  "000000001100010001",  "000000001100001100",  "000000001100000111",  "000000001100000011",  "000000001011111110",  "000000001011111001",  "000000001011110100",  "000000001011110000",  "000000001011101011",  "000000001011100110",  "000000001011100001",  "000000001011011101",  "000000001011011000",  "000000001011010011",  "000000001011001110",  "000000001011001010",  "000000001011000101",  "000000001011000000",  "000000001010111011",  "000000001010110110",  "000000001010110001",  "000000001010101101",  "000000001010101000",  "000000001010100011",  "000000001010011110",  "000000001010011001",  "000000001010010100",  "000000001010010000",  "000000001010001011",  "000000001010000110",  "000000001010000001",  "000000001001111100",  "000000001001110111",  "000000001001110010",  "000000001001101110",  "000000001001101001",  "000000001001100100",  "000000001001011111",  "000000001001011010",  "000000001001010101",  "000000001001010000",  "000000001001001011",  "000000001001000110",  "000000001001000001",  "000000001000111101",  "000000001000111000",  "000000001000110011",  "000000001000101110",  "000000001000101001",  "000000001000100100",  "000000001000011111",  "000000001000011010",  "000000001000010101",  "000000001000010000",  "000000001000001011",  "000000001000000110",  "000000001000000001",  "000000000111111100",  "000000000111110111",  "000000000111110010",  "000000000111101101",  "000000000111101000",  "000000000111100011",  "000000000111011111",  "000000000111011010",  "000000000111010101",  "000000000111010000",  "000000000111001011",  "000000000111000110",  "000000000111000001",  "000000000110111100",  "000000000110110111",  "000000000110110010",  "000000000110101101",  "000000000110101000",  "000000000110100011",  "000000000110011110",  "000000000110011001",  "000000000110010100",  "000000000110001111",  "000000000110001001",  "000000000110000100",  "000000000101111111",  "000000000101111010",  "000000000101110101",  "000000000101110000",  "000000000101101011",  "000000000101100110",  "000000000101100001",  "000000000101011100",  "000000000101010111",  "000000000101010010",  "000000000101001101",  "000000000101001000",  "000000000101000011",  "000000000100111110",  "000000000100111001",  "000000000100110100",  "000000000100101111",  "000000000100101010",  "000000000100100101",  "000000000100100000",  "000000000100011011",  "000000000100010110",  "000000000100010001",  "000000000100001100",  "000000000100000110",  "000000000100000001",  "000000000011111100",  "000000000011110111",  "000000000011110010",  "000000000011101101",  "000000000011101000",  "000000000011100011",  "000000000011011110",  "000000000011011001",  "000000000011010100",  "000000000011001111",  "000000000011001010",  "000000000011000101",  "000000000011000000",  "000000000010111011",  "000000000010110110",  "000000000010110001",  "000000000010101011",  "000000000010100110",  "000000000010100001",  "000000000010011100",  "000000000010010111",  "000000000010010010",  "000000000010001101",  "000000000010001000",  "000000000010000011",  "000000000001111110",  "000000000001111001",  "000000000001110100",  "000000000001101111",  "000000000001101010",  "000000000001100101",  "000000000001100000",  "000000000001011011",  "000000000001010110",  "000000000001010001",  "000000000001001100",  "000000000001000110",  "000000000001000001",  "000000000000111100",  "000000000000110111",  "000000000000110010",  "000000000000101101",  "000000000000101000",  "000000000000100011",  "000000000000011110",  "000000000000011001",  "000000000000010100",  "000000000000001111",  "000000000000001010",  "000000000000000101"),("000000000000000000",  "111111111111111011",  "111111111111110110",  "111111111111110001",  "111111111111101100",  "111111111111100111",  "111111111111100010",  "111111111111011101",  "111111111111011000",  "111111111111010011",  "111111111111001110",  "111111111111001001",  "111111111111000100",  "111111111110111111",  "111111111110111010",  "111111111110110101",  "111111111110110000",  "111111111110101011",  "111111111110100110",  "111111111110100001",  "111111111110011100",  "111111111110010111",  "111111111110010010",  "111111111110001101",  "111111111110001000",  "111111111110000011",  "111111111101111110",  "111111111101111001",  "111111111101110100",  "111111111101101111",  "111111111101101010",  "111111111101100101",  "111111111101100000",  "111111111101011100",  "111111111101010111",  "111111111101010010",  "111111111101001101",  "111111111101001000",  "111111111101000011",  "111111111100111110",  "111111111100111001",  "111111111100110100",  "111111111100101111",  "111111111100101010",  "111111111100100101",  "111111111100100001",  "111111111100011100",  "111111111100010111",  "111111111100010010",  "111111111100001101",  "111111111100001000",  "111111111100000011",  "111111111011111110",  "111111111011111010",  "111111111011110101",  "111111111011110000",  "111111111011101011",  "111111111011100110",  "111111111011100001",  "111111111011011100",  "111111111011011000",  "111111111011010011",  "111111111011001110",  "111111111011001001",  "111111111011000100",  "111111111011000000",  "111111111010111011",  "111111111010110110",  "111111111010110001",  "111111111010101100",  "111111111010101000",  "111111111010100011",  "111111111010011110",  "111111111010011001",  "111111111010010100",  "111111111010010000",  "111111111010001011",  "111111111010000110",  "111111111010000001",  "111111111001111101",  "111111111001111000",  "111111111001110011",  "111111111001101111",  "111111111001101010",  "111111111001100101",  "111111111001100000",  "111111111001011100",  "111111111001010111",  "111111111001010010",  "111111111001001110",  "111111111001001001",  "111111111001000100",  "111111111001000000",  "111111111000111011",  "111111111000110110",  "111111111000110010",  "111111111000101101",  "111111111000101000",  "111111111000100100",  "111111111000011111",  "111111111000011011",  "111111111000010110",  "111111111000010001",  "111111111000001101",  "111111111000001000",  "111111111000000100",  "111111110111111111",  "111111110111111010",  "111111110111110110",  "111111110111110001",  "111111110111101101",  "111111110111101000",  "111111110111100100",  "111111110111011111",  "111111110111011011",  "111111110111010110",  "111111110111010010",  "111111110111001101",  "111111110111001001",  "111111110111000100",  "111111110111000000",  "111111110110111011",  "111111110110110111",  "111111110110110010",  "111111110110101110",  "111111110110101001",  "111111110110100101",  "111111110110100000",  "111111110110011100",  "111111110110011000",  "111111110110010011",  "111111110110001111",  "111111110110001010",  "111111110110000110",  "111111110110000010",  "111111110101111101",  "111111110101111001",  "111111110101110100",  "111111110101110000",  "111111110101101100",  "111111110101100111",  "111111110101100011",  "111111110101011111",  "111111110101011010",  "111111110101010110",  "111111110101010010",  "111111110101001110",  "111111110101001001",  "111111110101000101",  "111111110101000001",  "111111110100111101",  "111111110100111000",  "111111110100110100",  "111111110100110000",  "111111110100101100",  "111111110100100111",  "111111110100100011",  "111111110100011111",  "111111110100011011",  "111111110100010111",  "111111110100010010",  "111111110100001110",  "111111110100001010",  "111111110100000110",  "111111110100000010",  "111111110011111110",  "111111110011111010",  "111111110011110101",  "111111110011110001",  "111111110011101101",  "111111110011101001",  "111111110011100101",  "111111110011100001",  "111111110011011101",  "111111110011011001",  "111111110011010101",  "111111110011010001",  "111111110011001101",  "111111110011001001",  "111111110011000101",  "111111110011000001",  "111111110010111101",  "111111110010111001",  "111111110010110101",  "111111110010110001",  "111111110010101101",  "111111110010101001",  "111111110010100101",  "111111110010100001",  "111111110010011101",  "111111110010011001",  "111111110010010110",  "111111110010010010",  "111111110010001110",  "111111110010001010",  "111111110010000110",  "111111110010000010",  "111111110001111110",  "111111110001111011",  "111111110001110111",  "111111110001110011",  "111111110001101111",  "111111110001101011",  "111111110001101000",  "111111110001100100",  "111111110001100000",  "111111110001011100",  "111111110001011001",  "111111110001010101",  "111111110001010001",  "111111110001001110",  "111111110001001010",  "111111110001000110",  "111111110001000011",  "111111110000111111",  "111111110000111011",  "111111110000111000",  "111111110000110100",  "111111110000110000",  "111111110000101101",  "111111110000101001",  "111111110000100110",  "111111110000100010",  "111111110000011110",  "111111110000011011",  "111111110000010111",  "111111110000010100",  "111111110000010000",  "111111110000001101",  "111111110000001001",  "111111110000000110",  "111111110000000010",  "111111101111111111",  "111111101111111011",  "111111101111111000",  "111111101111110101",  "111111101111110001",  "111111101111101110",  "111111101111101010",  "111111101111100111",  "111111101111100100",  "111111101111100000",  "111111101111011101",  "111111101111011001",  "111111101111010110",  "111111101111010011",  "111111101111010000",  "111111101111001100",  "111111101111001001",  "111111101111000110",  "111111101111000010",  "111111101110111111",  "111111101110111100",  "111111101110111001",  "111111101110110101",  "111111101110110010",  "111111101110101111",  "111111101110101100",  "111111101110101001",  "111111101110100110",  "111111101110100010",  "111111101110011111",  "111111101110011100",  "111111101110011001",  "111111101110010110",  "111111101110010011",  "111111101110010000",  "111111101110001101",  "111111101110001010",  "111111101110000111",  "111111101110000100",  "111111101110000001",  "111111101101111110",  "111111101101111011",  "111111101101111000",  "111111101101110101",  "111111101101110010",  "111111101101101111",  "111111101101101100",  "111111101101101001",  "111111101101100110",  "111111101101100011",  "111111101101100000",  "111111101101011101",  "111111101101011010",  "111111101101011000",  "111111101101010101",  "111111101101010010",  "111111101101001111",  "111111101101001100",  "111111101101001001",  "111111101101000111",  "111111101101000100",  "111111101101000001",  "111111101100111110",  "111111101100111100",  "111111101100111001",  "111111101100110110",  "111111101100110100",  "111111101100110001",  "111111101100101110",  "111111101100101100",  "111111101100101001",  "111111101100100110",  "111111101100100100",  "111111101100100001",  "111111101100011111",  "111111101100011100",  "111111101100011001",  "111111101100010111",  "111111101100010100",  "111111101100010010",  "111111101100001111",  "111111101100001101",  "111111101100001010",  "111111101100001000",  "111111101100000101",  "111111101100000011",  "111111101100000001",  "111111101011111110",  "111111101011111100",  "111111101011111001",  "111111101011110111",  "111111101011110101",  "111111101011110010",  "111111101011110000",  "111111101011101110",  "111111101011101011",  "111111101011101001",  "111111101011100111",  "111111101011100100",  "111111101011100010",  "111111101011100000",  "111111101011011110",  "111111101011011011",  "111111101011011001",  "111111101011010111",  "111111101011010101",  "111111101011010011",  "111111101011010001",  "111111101011001110",  "111111101011001100",  "111111101011001010",  "111111101011001000",  "111111101011000110",  "111111101011000100",  "111111101011000010",  "111111101011000000",  "111111101010111110",  "111111101010111100",  "111111101010111010",  "111111101010111000",  "111111101010110110",  "111111101010110100",  "111111101010110010",  "111111101010110000",  "111111101010101110",  "111111101010101100",  "111111101010101010",  "111111101010101000",  "111111101010100110",  "111111101010100101",  "111111101010100011",  "111111101010100001",  "111111101010011111",  "111111101010011101",  "111111101010011011",  "111111101010011010",  "111111101010011000",  "111111101010010110",  "111111101010010100",  "111111101010010011",  "111111101010010001",  "111111101010001111",  "111111101010001110",  "111111101010001100",  "111111101010001010",  "111111101010001001",  "111111101010000111",  "111111101010000101",  "111111101010000100",  "111111101010000010",  "111111101010000001",  "111111101001111111",  "111111101001111110",  "111111101001111100",  "111111101001111011",  "111111101001111001",  "111111101001111000",  "111111101001110110",  "111111101001110101",  "111111101001110011",  "111111101001110010",  "111111101001110000",  "111111101001101111",  "111111101001101110",  "111111101001101100",  "111111101001101011",  "111111101001101001",  "111111101001101000",  "111111101001100111",  "111111101001100110",  "111111101001100100",  "111111101001100011",  "111111101001100010",  "111111101001100000",  "111111101001011111",  "111111101001011110",  "111111101001011101",  "111111101001011100",  "111111101001011010",  "111111101001011001",  "111111101001011000",  "111111101001010111",  "111111101001010110",  "111111101001010101",  "111111101001010100",  "111111101001010011",  "111111101001010001",  "111111101001010000",  "111111101001001111",  "111111101001001110",  "111111101001001101",  "111111101001001100",  "111111101001001011",  "111111101001001010",  "111111101001001001",  "111111101001001001",  "111111101001001000",  "111111101001000111",  "111111101001000110",  "111111101001000101",  "111111101001000100",  "111111101001000011",  "111111101001000010",  "111111101001000010",  "111111101001000001",  "111111101001000000",  "111111101000111111",  "111111101000111110",  "111111101000111110",  "111111101000111101",  "111111101000111100",  "111111101000111011",  "111111101000111011",  "111111101000111010",  "111111101000111001",  "111111101000111001",  "111111101000111000",  "111111101000110111",  "111111101000110111",  "111111101000110110",  "111111101000110110",  "111111101000110101",  "111111101000110101",  "111111101000110100",  "111111101000110011",  "111111101000110011",  "111111101000110010",  "111111101000110010",  "111111101000110010",  "111111101000110001",  "111111101000110001",  "111111101000110000",  "111111101000110000",  "111111101000101111",  "111111101000101111",  "111111101000101111",  "111111101000101110",  "111111101000101110",  "111111101000101110",  "111111101000101101",  "111111101000101101",  "111111101000101101",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101010",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101011",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101100",  "111111101000101101",  "111111101000101101",  "111111101000101101",  "111111101000101110",  "111111101000101110",  "111111101000101110",  "111111101000101111",  "111111101000101111",  "111111101000101111",  "111111101000110000",  "111111101000110000",  "111111101000110001",  "111111101000110001",  "111111101000110001",  "111111101000110010",  "111111101000110010",  "111111101000110011",  "111111101000110011",  "111111101000110100",  "111111101000110100",  "111111101000110101",  "111111101000110101",  "111111101000110110",  "111111101000110111",  "111111101000110111",  "111111101000111000",  "111111101000111000",  "111111101000111001",  "111111101000111010",  "111111101000111010",  "111111101000111011",  "111111101000111100",  "111111101000111101",  "111111101000111101",  "111111101000111110",  "111111101000111111",  "111111101000111111",  "111111101001000000",  "111111101001000001",  "111111101001000010",  "111111101001000011",  "111111101001000100",  "111111101001000100",  "111111101001000101",  "111111101001000110",  "111111101001000111",  "111111101001001000",  "111111101001001001",  "111111101001001010",  "111111101001001011",  "111111101001001100",  "111111101001001101",  "111111101001001110",  "111111101001001111",  "111111101001010000",  "111111101001010001",  "111111101001010010",  "111111101001010011",  "111111101001010100",  "111111101001010101",  "111111101001010110",  "111111101001010111",  "111111101001011000",  "111111101001011001",  "111111101001011010",  "111111101001011100",  "111111101001011101",  "111111101001011110",  "111111101001011111",  "111111101001100000",  "111111101001100001",  "111111101001100011",  "111111101001100100",  "111111101001100101",  "111111101001100110",  "111111101001101000",  "111111101001101001",  "111111101001101010",  "111111101001101100",  "111111101001101101",  "111111101001101110",  "111111101001110000",  "111111101001110001",  "111111101001110011",  "111111101001110100",  "111111101001110101",  "111111101001110111",  "111111101001111000",  "111111101001111010",  "111111101001111011",  "111111101001111101",  "111111101001111110",  "111111101010000000",  "111111101010000001",  "111111101010000011",  "111111101010000100",  "111111101010000110",  "111111101010000111",  "111111101010001001",  "111111101010001010",  "111111101010001100",  "111111101010001110",  "111111101010001111",  "111111101010010001",  "111111101010010011",  "111111101010010100",  "111111101010010110",  "111111101010011000",  "111111101010011001",  "111111101010011011",  "111111101010011101",  "111111101010011111",  "111111101010100000",  "111111101010100010",  "111111101010100100",  "111111101010100110",  "111111101010101000",  "111111101010101001",  "111111101010101011",  "111111101010101101",  "111111101010101111",  "111111101010110001",  "111111101010110011",  "111111101010110100",  "111111101010110110",  "111111101010111000",  "111111101010111010",  "111111101010111100",  "111111101010111110",  "111111101011000000",  "111111101011000010",  "111111101011000100",  "111111101011000110",  "111111101011001000",  "111111101011001010",  "111111101011001100",  "111111101011001110",  "111111101011010000",  "111111101011010010",  "111111101011010100",  "111111101011010110",  "111111101011011001",  "111111101011011011",  "111111101011011101",  "111111101011011111",  "111111101011100001",  "111111101011100011",  "111111101011100101",  "111111101011101000",  "111111101011101010",  "111111101011101100",  "111111101011101110",  "111111101011110001",  "111111101011110011",  "111111101011110101",  "111111101011110111",  "111111101011111010",  "111111101011111100",  "111111101011111110",  "111111101100000000",  "111111101100000011",  "111111101100000101",  "111111101100000111",  "111111101100001010",  "111111101100001100",  "111111101100001111",  "111111101100010001",  "111111101100010011",  "111111101100010110",  "111111101100011000",  "111111101100011011",  "111111101100011101",  "111111101100100000",  "111111101100100010",  "111111101100100100",  "111111101100100111",  "111111101100101001",  "111111101100101100",  "111111101100101110",  "111111101100110001",  "111111101100110100",  "111111101100110110",  "111111101100111001",  "111111101100111011",  "111111101100111110",  "111111101101000000",  "111111101101000011",  "111111101101000110",  "111111101101001000",  "111111101101001011",  "111111101101001110",  "111111101101010000",  "111111101101010011",  "111111101101010110",  "111111101101011000",  "111111101101011011",  "111111101101011110",  "111111101101100000",  "111111101101100011",  "111111101101100110",  "111111101101101001",  "111111101101101011",  "111111101101101110",  "111111101101110001",  "111111101101110100",  "111111101101110111",  "111111101101111001",  "111111101101111100",  "111111101101111111",  "111111101110000010",  "111111101110000101",  "111111101110001000",  "111111101110001010",  "111111101110001101",  "111111101110010000",  "111111101110010011",  "111111101110010110",  "111111101110011001",  "111111101110011100",  "111111101110011111",  "111111101110100010",  "111111101110100101",  "111111101110101000",  "111111101110101011",  "111111101110101110",  "111111101110110001",  "111111101110110100",  "111111101110110111",  "111111101110111010",  "111111101110111101",  "111111101111000000",  "111111101111000011",  "111111101111000110",  "111111101111001001",  "111111101111001100",  "111111101111001111",  "111111101111010010",  "111111101111010101",  "111111101111011000",  "111111101111011011",  "111111101111011111",  "111111101111100010",  "111111101111100101",  "111111101111101000",  "111111101111101011",  "111111101111101110",  "111111101111110010",  "111111101111110101",  "111111101111111000",  "111111101111111011",  "111111101111111110",  "111111110000000010",  "111111110000000101",  "111111110000001000",  "111111110000001011",  "111111110000001111",  "111111110000010010",  "111111110000010101",  "111111110000011000",  "111111110000011100",  "111111110000011111",  "111111110000100010",  "111111110000100110",  "111111110000101001",  "111111110000101100",  "111111110000110000",  "111111110000110011",  "111111110000110110",  "111111110000111010",  "111111110000111101",  "111111110001000000",  "111111110001000100",  "111111110001000111",  "111111110001001011",  "111111110001001110",  "111111110001010001",  "111111110001010101",  "111111110001011000",  "111111110001011100",  "111111110001011111",  "111111110001100011",  "111111110001100110",  "111111110001101010",  "111111110001101101",  "111111110001110001",  "111111110001110100",  "111111110001111000",  "111111110001111011",  "111111110001111111",  "111111110010000010",  "111111110010000110",  "111111110010001001",  "111111110010001101",  "111111110010010000",  "111111110010010100",  "111111110010010111",  "111111110010011011",  "111111110010011111",  "111111110010100010",  "111111110010100110",  "111111110010101001",  "111111110010101101",  "111111110010110001",  "111111110010110100",  "111111110010111000",  "111111110010111011",  "111111110010111111",  "111111110011000011",  "111111110011000110",  "111111110011001010",  "111111110011001110",  "111111110011010001",  "111111110011010101",  "111111110011011001",  "111111110011011100",  "111111110011100000",  "111111110011100100",  "111111110011101000",  "111111110011101011",  "111111110011101111",  "111111110011110011",  "111111110011110110",  "111111110011111010",  "111111110011111110",  "111111110100000010",  "111111110100000101",  "111111110100001001",  "111111110100001101",  "111111110100010001",  "111111110100010101",  "111111110100011000",  "111111110100011100",  "111111110100100000",  "111111110100100100",  "111111110100101000",  "111111110100101011",  "111111110100101111",  "111111110100110011",  "111111110100110111",  "111111110100111011",  "111111110100111111",  "111111110101000010",  "111111110101000110",  "111111110101001010",  "111111110101001110",  "111111110101010010",  "111111110101010110",  "111111110101011010",  "111111110101011101",  "111111110101100001",  "111111110101100101",  "111111110101101001",  "111111110101101101",  "111111110101110001",  "111111110101110101",  "111111110101111001",  "111111110101111101",  "111111110110000001",  "111111110110000101",  "111111110110001000",  "111111110110001100",  "111111110110010000",  "111111110110010100",  "111111110110011000",  "111111110110011100",  "111111110110100000",  "111111110110100100",  "111111110110101000",  "111111110110101100",  "111111110110110000",  "111111110110110100",  "111111110110111000",  "111111110110111100",  "111111110111000000",  "111111110111000100",  "111111110111001000",  "111111110111001100",  "111111110111010000",  "111111110111010100",  "111111110111011000",  "111111110111011100",  "111111110111100000",  "111111110111100100",  "111111110111101000",  "111111110111101100",  "111111110111110000",  "111111110111110100",  "111111110111111000",  "111111110111111100",  "111111111000000000",  "111111111000000100",  "111111111000001001",  "111111111000001101",  "111111111000010001",  "111111111000010101",  "111111111000011001",  "111111111000011101",  "111111111000100001",  "111111111000100101",  "111111111000101001",  "111111111000101101",  "111111111000110001",  "111111111000110101",  "111111111000111001",  "111111111000111110",  "111111111001000010",  "111111111001000110",  "111111111001001010",  "111111111001001110",  "111111111001010010",  "111111111001010110",  "111111111001011010",  "111111111001011110",  "111111111001100011",  "111111111001100111",  "111111111001101011",  "111111111001101111",  "111111111001110011",  "111111111001110111",  "111111111001111011",  "111111111010000000",  "111111111010000100",  "111111111010001000",  "111111111010001100",  "111111111010010000",  "111111111010010100",  "111111111010011000",  "111111111010011101",  "111111111010100001",  "111111111010100101",  "111111111010101001",  "111111111010101101",  "111111111010110001",  "111111111010110101",  "111111111010111010",  "111111111010111110",  "111111111011000010",  "111111111011000110",  "111111111011001010",  "111111111011001110",  "111111111011010011",  "111111111011010111",  "111111111011011011",  "111111111011011111",  "111111111011100011",  "111111111011101000",  "111111111011101100",  "111111111011110000",  "111111111011110100",  "111111111011111000",  "111111111011111100",  "111111111100000001",  "111111111100000101",  "111111111100001001",  "111111111100001101",  "111111111100010001",  "111111111100010110",  "111111111100011010",  "111111111100011110",  "111111111100100010",  "111111111100100110",  "111111111100101011",  "111111111100101111",  "111111111100110011",  "111111111100110111",  "111111111100111011",  "111111111100111111",  "111111111101000100",  "111111111101001000",  "111111111101001100",  "111111111101010000",  "111111111101010100",  "111111111101011001",  "111111111101011101",  "111111111101100001",  "111111111101100101",  "111111111101101001",  "111111111101101110",  "111111111101110010",  "111111111101110110",  "111111111101111010",  "111111111101111110",  "111111111110000011",  "111111111110000111",  "111111111110001011",  "111111111110001111",  "111111111110010011",  "111111111110011000",  "111111111110011100",  "111111111110100000",  "111111111110100100",  "111111111110101000",  "111111111110101100",  "111111111110110001",  "111111111110110101",  "111111111110111001",  "111111111110111101",  "111111111111000001",  "111111111111000110",  "111111111111001010",  "111111111111001110",  "111111111111010010",  "111111111111010110",  "111111111111011010",  "111111111111011111",  "111111111111100011",  "111111111111100111",  "111111111111101011",  "111111111111101111",  "111111111111110100",  "111111111111111000",  "111111111111111100"),("000000000000000000",  "000000000000000100",  "000000000000001000",  "000000000000001100",  "000000000000010001",  "000000000000010101",  "000000000000011001",  "000000000000011101",  "000000000000100001",  "000000000000100101",  "000000000000101010",  "000000000000101110",  "000000000000110010",  "000000000000110110",  "000000000000111010",  "000000000000111110",  "000000000001000010",  "000000000001000111",  "000000000001001011",  "000000000001001111",  "000000000001010011",  "000000000001010111",  "000000000001011011",  "000000000001011111",  "000000000001100011",  "000000000001101000",  "000000000001101100",  "000000000001110000",  "000000000001110100",  "000000000001111000",  "000000000001111100",  "000000000010000000",  "000000000010000100",  "000000000010001000",  "000000000010001100",  "000000000010010001",  "000000000010010101",  "000000000010011001",  "000000000010011101",  "000000000010100001",  "000000000010100101",  "000000000010101001",  "000000000010101101",  "000000000010110001",  "000000000010110101",  "000000000010111001",  "000000000010111101",  "000000000011000001",  "000000000011000101",  "000000000011001001",  "000000000011001101",  "000000000011010001",  "000000000011010110",  "000000000011011010",  "000000000011011110",  "000000000011100010",  "000000000011100110",  "000000000011101010",  "000000000011101110",  "000000000011110010",  "000000000011110110",  "000000000011111010",  "000000000011111110",  "000000000100000010",  "000000000100000110",  "000000000100001010",  "000000000100001110",  "000000000100010010",  "000000000100010110",  "000000000100011010",  "000000000100011101",  "000000000100100001",  "000000000100100101",  "000000000100101001",  "000000000100101101",  "000000000100110001",  "000000000100110101",  "000000000100111001",  "000000000100111101",  "000000000101000001",  "000000000101000101",  "000000000101001001",  "000000000101001101",  "000000000101010001",  "000000000101010101",  "000000000101011000",  "000000000101011100",  "000000000101100000",  "000000000101100100",  "000000000101101000",  "000000000101101100",  "000000000101110000",  "000000000101110100",  "000000000101110111",  "000000000101111011",  "000000000101111111",  "000000000110000011",  "000000000110000111",  "000000000110001011",  "000000000110001111",  "000000000110010010",  "000000000110010110",  "000000000110011010",  "000000000110011110",  "000000000110100010",  "000000000110100101",  "000000000110101001",  "000000000110101101",  "000000000110110001",  "000000000110110101",  "000000000110111000",  "000000000110111100",  "000000000111000000",  "000000000111000100",  "000000000111000111",  "000000000111001011",  "000000000111001111",  "000000000111010011",  "000000000111010110",  "000000000111011010",  "000000000111011110",  "000000000111100001",  "000000000111100101",  "000000000111101001",  "000000000111101100",  "000000000111110000",  "000000000111110100",  "000000000111110111",  "000000000111111011",  "000000000111111111",  "000000001000000010",  "000000001000000110",  "000000001000001010",  "000000001000001101",  "000000001000010001",  "000000001000010101",  "000000001000011000",  "000000001000011100",  "000000001000011111",  "000000001000100011",  "000000001000100111",  "000000001000101010",  "000000001000101110",  "000000001000110001",  "000000001000110101",  "000000001000111001",  "000000001000111100",  "000000001001000000",  "000000001001000011",  "000000001001000111",  "000000001001001010",  "000000001001001110",  "000000001001010001",  "000000001001010101",  "000000001001011000",  "000000001001011100",  "000000001001011111",  "000000001001100011",  "000000001001100110",  "000000001001101010",  "000000001001101101",  "000000001001110000",  "000000001001110100",  "000000001001110111",  "000000001001111011",  "000000001001111110",  "000000001010000010",  "000000001010000101",  "000000001010001000",  "000000001010001100",  "000000001010001111",  "000000001010010011",  "000000001010010110",  "000000001010011001",  "000000001010011101",  "000000001010100000",  "000000001010100011",  "000000001010100111",  "000000001010101010",  "000000001010101101",  "000000001010110001",  "000000001010110100",  "000000001010110111",  "000000001010111010",  "000000001010111110",  "000000001011000001",  "000000001011000100",  "000000001011000111",  "000000001011001011",  "000000001011001110",  "000000001011010001",  "000000001011010100",  "000000001011011000",  "000000001011011011",  "000000001011011110",  "000000001011100001",  "000000001011100100",  "000000001011100111",  "000000001011101011",  "000000001011101110",  "000000001011110001",  "000000001011110100",  "000000001011110111",  "000000001011111010",  "000000001011111101",  "000000001100000001",  "000000001100000100",  "000000001100000111",  "000000001100001010",  "000000001100001101",  "000000001100010000",  "000000001100010011",  "000000001100010110",  "000000001100011001",  "000000001100011100",  "000000001100011111",  "000000001100100010",  "000000001100100101",  "000000001100101000",  "000000001100101011",  "000000001100101110",  "000000001100110001",  "000000001100110100",  "000000001100110111",  "000000001100111010",  "000000001100111101",  "000000001101000000",  "000000001101000011",  "000000001101000110",  "000000001101001000",  "000000001101001011",  "000000001101001110",  "000000001101010001",  "000000001101010100",  "000000001101010111",  "000000001101011010",  "000000001101011100",  "000000001101011111",  "000000001101100010",  "000000001101100101",  "000000001101101000",  "000000001101101010",  "000000001101101101",  "000000001101110000",  "000000001101110011",  "000000001101110101",  "000000001101111000",  "000000001101111011",  "000000001101111110",  "000000001110000000",  "000000001110000011",  "000000001110000110",  "000000001110001000",  "000000001110001011",  "000000001110001110",  "000000001110010000",  "000000001110010011",  "000000001110010110",  "000000001110011000",  "000000001110011011",  "000000001110011101",  "000000001110100000",  "000000001110100011",  "000000001110100101",  "000000001110101000",  "000000001110101010",  "000000001110101101",  "000000001110101111",  "000000001110110010",  "000000001110110100",  "000000001110110111",  "000000001110111001",  "000000001110111100",  "000000001110111110",  "000000001111000001",  "000000001111000011",  "000000001111000110",  "000000001111001000",  "000000001111001011",  "000000001111001101",  "000000001111001111",  "000000001111010010",  "000000001111010100",  "000000001111010111",  "000000001111011001",  "000000001111011011",  "000000001111011110",  "000000001111100000",  "000000001111100010",  "000000001111100101",  "000000001111100111",  "000000001111101001",  "000000001111101100",  "000000001111101110",  "000000001111110000",  "000000001111110010",  "000000001111110101",  "000000001111110111",  "000000001111111001",  "000000001111111011",  "000000001111111101",  "000000010000000000",  "000000010000000010",  "000000010000000100",  "000000010000000110",  "000000010000001000",  "000000010000001010",  "000000010000001101",  "000000010000001111",  "000000010000010001",  "000000010000010011",  "000000010000010101",  "000000010000010111",  "000000010000011001",  "000000010000011011",  "000000010000011101",  "000000010000011111",  "000000010000100001",  "000000010000100011",  "000000010000100101",  "000000010000100111",  "000000010000101001",  "000000010000101011",  "000000010000101101",  "000000010000101111",  "000000010000110001",  "000000010000110011",  "000000010000110101",  "000000010000110111",  "000000010000111001",  "000000010000111010",  "000000010000111100",  "000000010000111110",  "000000010001000000",  "000000010001000010",  "000000010001000100",  "000000010001000101",  "000000010001000111",  "000000010001001001",  "000000010001001011",  "000000010001001101",  "000000010001001110",  "000000010001010000",  "000000010001010010",  "000000010001010100",  "000000010001010101",  "000000010001010111",  "000000010001011001",  "000000010001011010",  "000000010001011100",  "000000010001011110",  "000000010001011111",  "000000010001100001",  "000000010001100011",  "000000010001100100",  "000000010001100110",  "000000010001100111",  "000000010001101001",  "000000010001101011",  "000000010001101100",  "000000010001101110",  "000000010001101111",  "000000010001110001",  "000000010001110010",  "000000010001110100",  "000000010001110101",  "000000010001110111",  "000000010001111000",  "000000010001111010",  "000000010001111011",  "000000010001111100",  "000000010001111110",  "000000010001111111",  "000000010010000001",  "000000010010000010",  "000000010010000011",  "000000010010000101",  "000000010010000110",  "000000010010000111",  "000000010010001001",  "000000010010001010",  "000000010010001011",  "000000010010001101",  "000000010010001110",  "000000010010001111",  "000000010010010001",  "000000010010010010",  "000000010010010011",  "000000010010010100",  "000000010010010101",  "000000010010010111",  "000000010010011000",  "000000010010011001",  "000000010010011010",  "000000010010011011",  "000000010010011100",  "000000010010011110",  "000000010010011111",  "000000010010100000",  "000000010010100001",  "000000010010100010",  "000000010010100011",  "000000010010100100",  "000000010010100101",  "000000010010100110",  "000000010010100111",  "000000010010101000",  "000000010010101001",  "000000010010101010",  "000000010010101011",  "000000010010101100",  "000000010010101101",  "000000010010101110",  "000000010010101111",  "000000010010110000",  "000000010010110001",  "000000010010110010",  "000000010010110011",  "000000010010110100",  "000000010010110100",  "000000010010110101",  "000000010010110110",  "000000010010110111",  "000000010010111000",  "000000010010111001",  "000000010010111001",  "000000010010111010",  "000000010010111011",  "000000010010111100",  "000000010010111100",  "000000010010111101",  "000000010010111110",  "000000010010111111",  "000000010010111111",  "000000010011000000",  "000000010011000001",  "000000010011000001",  "000000010011000010",  "000000010011000011",  "000000010011000011",  "000000010011000100",  "000000010011000100",  "000000010011000101",  "000000010011000110",  "000000010011000110",  "000000010011000111",  "000000010011000111",  "000000010011001000",  "000000010011001000",  "000000010011001001",  "000000010011001001",  "000000010011001010",  "000000010011001010",  "000000010011001011",  "000000010011001011",  "000000010011001100",  "000000010011001100",  "000000010011001101",  "000000010011001101",  "000000010011001101",  "000000010011001110",  "000000010011001110",  "000000010011001110",  "000000010011001111",  "000000010011001111",  "000000010011001111",  "000000010011010000",  "000000010011010000",  "000000010011010000",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010100",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010011",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010010",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010001",  "000000010011010000",  "000000010011010000",  "000000010011010000",  "000000010011010000",  "000000010011001111",  "000000010011001111",  "000000010011001111",  "000000010011001110",  "000000010011001110",  "000000010011001101",  "000000010011001101",  "000000010011001101",  "000000010011001100",  "000000010011001100",  "000000010011001011",  "000000010011001011",  "000000010011001010",  "000000010011001010",  "000000010011001010",  "000000010011001001",  "000000010011001001",  "000000010011001000",  "000000010011001000",  "000000010011000111",  "000000010011000110",  "000000010011000110",  "000000010011000101",  "000000010011000101",  "000000010011000100",  "000000010011000100",  "000000010011000011",  "000000010011000010",  "000000010011000010",  "000000010011000001",  "000000010011000000",  "000000010011000000",  "000000010010111111",  "000000010010111110",  "000000010010111110",  "000000010010111101",  "000000010010111100",  "000000010010111011",  "000000010010111011",  "000000010010111010",  "000000010010111001",  "000000010010111000",  "000000010010111000",  "000000010010110111",  "000000010010110110",  "000000010010110101",  "000000010010110100",  "000000010010110011",  "000000010010110011",  "000000010010110010",  "000000010010110001",  "000000010010110000",  "000000010010101111",  "000000010010101110",  "000000010010101101",  "000000010010101100",  "000000010010101011",  "000000010010101010",  "000000010010101001",  "000000010010101000",  "000000010010100111",  "000000010010100110",  "000000010010100101",  "000000010010100100",  "000000010010100011",  "000000010010100010",  "000000010010100001",  "000000010010100000",  "000000010010011111",  "000000010010011110",  "000000010010011101",  "000000010010011100",  "000000010010011011",  "000000010010011001",  "000000010010011000",  "000000010010010111",  "000000010010010110",  "000000010010010101",  "000000010010010100",  "000000010010010010",  "000000010010010001",  "000000010010010000",  "000000010010001111",  "000000010010001110",  "000000010010001100",  "000000010010001011",  "000000010010001010",  "000000010010001000",  "000000010010000111",  "000000010010000110",  "000000010010000101",  "000000010010000011",  "000000010010000010",  "000000010010000001",  "000000010001111111",  "000000010001111110",  "000000010001111100",  "000000010001111011",  "000000010001111010",  "000000010001111000",  "000000010001110111",  "000000010001110101",  "000000010001110100",  "000000010001110011",  "000000010001110001",  "000000010001110000",  "000000010001101110",  "000000010001101101",  "000000010001101011",  "000000010001101010",  "000000010001101000",  "000000010001100111",  "000000010001100101",  "000000010001100100",  "000000010001100010",  "000000010001100000",  "000000010001011111",  "000000010001011101",  "000000010001011100",  "000000010001011010",  "000000010001011000",  "000000010001010111",  "000000010001010101",  "000000010001010011",  "000000010001010010",  "000000010001010000",  "000000010001001110",  "000000010001001101",  "000000010001001011",  "000000010001001001",  "000000010001001000",  "000000010001000110",  "000000010001000100",  "000000010001000010",  "000000010001000001",  "000000010000111111",  "000000010000111101",  "000000010000111011",  "000000010000111010",  "000000010000111000",  "000000010000110110",  "000000010000110100",  "000000010000110010",  "000000010000110000",  "000000010000101111",  "000000010000101101",  "000000010000101011",  "000000010000101001",  "000000010000100111",  "000000010000100101",  "000000010000100011",  "000000010000100001",  "000000010000011111",  "000000010000011110",  "000000010000011100",  "000000010000011010",  "000000010000011000",  "000000010000010110",  "000000010000010100",  "000000010000010010",  "000000010000010000",  "000000010000001110",  "000000010000001100",  "000000010000001010",  "000000010000001000",  "000000010000000110",  "000000010000000100",  "000000010000000001",  "000000001111111111",  "000000001111111101",  "000000001111111011",  "000000001111111001",  "000000001111110111",  "000000001111110101",  "000000001111110011",  "000000001111110001",  "000000001111101111",  "000000001111101100",  "000000001111101010",  "000000001111101000",  "000000001111100110",  "000000001111100100",  "000000001111100001",  "000000001111011111",  "000000001111011101",  "000000001111011011",  "000000001111011001",  "000000001111010110",  "000000001111010100",  "000000001111010010",  "000000001111010000",  "000000001111001101",  "000000001111001011",  "000000001111001001",  "000000001111000111",  "000000001111000100",  "000000001111000010",  "000000001111000000",  "000000001110111101",  "000000001110111011",  "000000001110111001",  "000000001110110110",  "000000001110110100",  "000000001110110001",  "000000001110101111",  "000000001110101101",  "000000001110101010",  "000000001110101000",  "000000001110100110",  "000000001110100011",  "000000001110100001",  "000000001110011110",  "000000001110011100",  "000000001110011001",  "000000001110010111",  "000000001110010100",  "000000001110010010",  "000000001110010000",  "000000001110001101",  "000000001110001011",  "000000001110001000",  "000000001110000110",  "000000001110000011",  "000000001110000000",  "000000001101111110",  "000000001101111011",  "000000001101111001",  "000000001101110110",  "000000001101110100",  "000000001101110001",  "000000001101101111",  "000000001101101100",  "000000001101101001",  "000000001101100111",  "000000001101100100",  "000000001101100010",  "000000001101011111",  "000000001101011100",  "000000001101011010",  "000000001101010111",  "000000001101010100",  "000000001101010010",  "000000001101001111",  "000000001101001100",  "000000001101001010",  "000000001101000111",  "000000001101000100",  "000000001101000010",  "000000001100111111",  "000000001100111100",  "000000001100111010",  "000000001100110111",  "000000001100110100",  "000000001100110001",  "000000001100101111",  "000000001100101100",  "000000001100101001",  "000000001100100110",  "000000001100100100",  "000000001100100001",  "000000001100011110",  "000000001100011011",  "000000001100011000",  "000000001100010110",  "000000001100010011",  "000000001100010000",  "000000001100001101",  "000000001100001010",  "000000001100001000",  "000000001100000101",  "000000001100000010",  "000000001011111111",  "000000001011111100",  "000000001011111001",  "000000001011110110",  "000000001011110100",  "000000001011110001",  "000000001011101110",  "000000001011101011",  "000000001011101000",  "000000001011100101",  "000000001011100010",  "000000001011011111",  "000000001011011100",  "000000001011011001",  "000000001011010110",  "000000001011010011",  "000000001011010001",  "000000001011001110",  "000000001011001011",  "000000001011001000",  "000000001011000101",  "000000001011000010",  "000000001010111111",  "000000001010111100",  "000000001010111001",  "000000001010110110",  "000000001010110011",  "000000001010110000",  "000000001010101101",  "000000001010101010",  "000000001010100111",  "000000001010100100",  "000000001010100001",  "000000001010011110",  "000000001010011011",  "000000001010010111",  "000000001010010100",  "000000001010010001",  "000000001010001110",  "000000001010001011",  "000000001010001000",  "000000001010000101",  "000000001010000010",  "000000001001111111",  "000000001001111100",  "000000001001111001",  "000000001001110110",  "000000001001110010",  "000000001001101111",  "000000001001101100",  "000000001001101001",  "000000001001100110",  "000000001001100011",  "000000001001100000",  "000000001001011101",  "000000001001011001",  "000000001001010110",  "000000001001010011",  "000000001001010000",  "000000001001001101",  "000000001001001010",  "000000001001000110",  "000000001001000011",  "000000001001000000",  "000000001000111101",  "000000001000111010",  "000000001000110110",  "000000001000110011",  "000000001000110000",  "000000001000101101",  "000000001000101010",  "000000001000100110",  "000000001000100011",  "000000001000100000",  "000000001000011101",  "000000001000011010",  "000000001000010110",  "000000001000010011",  "000000001000010000",  "000000001000001101",  "000000001000001001",  "000000001000000110",  "000000001000000011",  "000000001000000000",  "000000000111111100",  "000000000111111001",  "000000000111110110",  "000000000111110010",  "000000000111101111",  "000000000111101100",  "000000000111101001",  "000000000111100101",  "000000000111100010",  "000000000111011111",  "000000000111011011",  "000000000111011000",  "000000000111010101",  "000000000111010010",  "000000000111001110",  "000000000111001011",  "000000000111001000",  "000000000111000100",  "000000000111000001",  "000000000110111110",  "000000000110111010",  "000000000110110111",  "000000000110110100",  "000000000110110000",  "000000000110101101",  "000000000110101010",  "000000000110100110",  "000000000110100011",  "000000000110100000",  "000000000110011100",  "000000000110011001",  "000000000110010101",  "000000000110010010",  "000000000110001111",  "000000000110001011",  "000000000110001000",  "000000000110000101",  "000000000110000001",  "000000000101111110",  "000000000101111010",  "000000000101110111",  "000000000101110100",  "000000000101110000",  "000000000101101101",  "000000000101101010",  "000000000101100110",  "000000000101100011",  "000000000101011111",  "000000000101011100",  "000000000101011001",  "000000000101010101",  "000000000101010010",  "000000000101001110",  "000000000101001011",  "000000000101001000",  "000000000101000100",  "000000000101000001",  "000000000100111101",  "000000000100111010",  "000000000100110110",  "000000000100110011",  "000000000100110000",  "000000000100101100",  "000000000100101001",  "000000000100100101",  "000000000100100010",  "000000000100011110",  "000000000100011011",  "000000000100011000",  "000000000100010100",  "000000000100010001",  "000000000100001101",  "000000000100001010",  "000000000100000110",  "000000000100000011",  "000000000100000000",  "000000000011111100",  "000000000011111001",  "000000000011110101",  "000000000011110010",  "000000000011101110",  "000000000011101011",  "000000000011100111",  "000000000011100100",  "000000000011100001",  "000000000011011101",  "000000000011011010",  "000000000011010110",  "000000000011010011",  "000000000011001111",  "000000000011001100",  "000000000011001000",  "000000000011000101",  "000000000011000001",  "000000000010111110",  "000000000010111011",  "000000000010110111",  "000000000010110100",  "000000000010110000",  "000000000010101101",  "000000000010101001",  "000000000010100110",  "000000000010100010",  "000000000010011111",  "000000000010011011",  "000000000010011000",  "000000000010010100",  "000000000010010001",  "000000000010001110",  "000000000010001010",  "000000000010000111",  "000000000010000011",  "000000000010000000",  "000000000001111100",  "000000000001111001",  "000000000001110101",  "000000000001110010",  "000000000001101110",  "000000000001101011",  "000000000001100111",  "000000000001100100",  "000000000001100001",  "000000000001011101",  "000000000001011010",  "000000000001010110",  "000000000001010011",  "000000000001001111",  "000000000001001100",  "000000000001001000",  "000000000001000101",  "000000000001000001",  "000000000000111110",  "000000000000111011",  "000000000000110111",  "000000000000110100",  "000000000000110000",  "000000000000101101",  "000000000000101001",  "000000000000100110",  "000000000000100010",  "000000000000011111",  "000000000000011100",  "000000000000011000",  "000000000000010101",  "000000000000010001",  "000000000000001110",  "000000000000001010",  "000000000000000111",  "000000000000000011"),("000000000000000000",  "111111111111111101",  "111111111111111001",  "111111111111110110",  "111111111111110010",  "111111111111101111",  "111111111111101011",  "111111111111101000",  "111111111111100101",  "111111111111100001",  "111111111111011110",  "111111111111011010",  "111111111111010111",  "111111111111010011",  "111111111111010000",  "111111111111001101",  "111111111111001001",  "111111111111000110",  "111111111111000010",  "111111111110111111",  "111111111110111100",  "111111111110111000",  "111111111110110101",  "111111111110110001",  "111111111110101110",  "111111111110101011",  "111111111110100111",  "111111111110100100",  "111111111110100000",  "111111111110011101",  "111111111110011010",  "111111111110010110",  "111111111110010011",  "111111111110010000",  "111111111110001100",  "111111111110001001",  "111111111110000101",  "111111111110000010",  "111111111101111111",  "111111111101111011",  "111111111101111000",  "111111111101110101",  "111111111101110001",  "111111111101101110",  "111111111101101011",  "111111111101100111",  "111111111101100100",  "111111111101100001",  "111111111101011101",  "111111111101011010",  "111111111101010111",  "111111111101010011",  "111111111101010000",  "111111111101001101",  "111111111101001001",  "111111111101000110",  "111111111101000011",  "111111111100111111",  "111111111100111100",  "111111111100111001",  "111111111100110101",  "111111111100110010",  "111111111100101111",  "111111111100101100",  "111111111100101000",  "111111111100100101",  "111111111100100010",  "111111111100011110",  "111111111100011011",  "111111111100011000",  "111111111100010101",  "111111111100010001",  "111111111100001110",  "111111111100001011",  "111111111100001000",  "111111111100000100",  "111111111100000001",  "111111111011111110",  "111111111011111011",  "111111111011110111",  "111111111011110100",  "111111111011110001",  "111111111011101110",  "111111111011101010",  "111111111011100111",  "111111111011100100",  "111111111011100001",  "111111111011011110",  "111111111011011010",  "111111111011010111",  "111111111011010100",  "111111111011010001",  "111111111011001110",  "111111111011001011",  "111111111011000111",  "111111111011000100",  "111111111011000001",  "111111111010111110",  "111111111010111011",  "111111111010111000",  "111111111010110100",  "111111111010110001",  "111111111010101110",  "111111111010101011",  "111111111010101000",  "111111111010100101",  "111111111010100010",  "111111111010011110",  "111111111010011011",  "111111111010011000",  "111111111010010101",  "111111111010010010",  "111111111010001111",  "111111111010001100",  "111111111010001001",  "111111111010000110",  "111111111010000011",  "111111111010000000",  "111111111001111100",  "111111111001111001",  "111111111001110110",  "111111111001110011",  "111111111001110000",  "111111111001101101",  "111111111001101010",  "111111111001100111",  "111111111001100100",  "111111111001100001",  "111111111001011110",  "111111111001011011",  "111111111001011000",  "111111111001010101",  "111111111001010010",  "111111111001001111",  "111111111001001100",  "111111111001001001",  "111111111001000110",  "111111111001000011",  "111111111001000000",  "111111111000111101",  "111111111000111010",  "111111111000110111",  "111111111000110100",  "111111111000110001",  "111111111000101110",  "111111111000101100",  "111111111000101001",  "111111111000100110",  "111111111000100011",  "111111111000100000",  "111111111000011101",  "111111111000011010",  "111111111000010111",  "111111111000010100",  "111111111000010001",  "111111111000001111",  "111111111000001100",  "111111111000001001",  "111111111000000110",  "111111111000000011",  "111111111000000000",  "111111110111111101",  "111111110111111011",  "111111110111111000",  "111111110111110101",  "111111110111110010",  "111111110111101111",  "111111110111101101",  "111111110111101010",  "111111110111100111",  "111111110111100100",  "111111110111100001",  "111111110111011111",  "111111110111011100",  "111111110111011001",  "111111110111010110",  "111111110111010100",  "111111110111010001",  "111111110111001110",  "111111110111001011",  "111111110111001001",  "111111110111000110",  "111111110111000011",  "111111110111000001",  "111111110110111110",  "111111110110111011",  "111111110110111001",  "111111110110110110",  "111111110110110011",  "111111110110110001",  "111111110110101110",  "111111110110101011",  "111111110110101001",  "111111110110100110",  "111111110110100011",  "111111110110100001",  "111111110110011110",  "111111110110011100",  "111111110110011001",  "111111110110010110",  "111111110110010100",  "111111110110010001",  "111111110110001111",  "111111110110001100",  "111111110110001001",  "111111110110000111",  "111111110110000100",  "111111110110000010",  "111111110101111111",  "111111110101111101",  "111111110101111010",  "111111110101111000",  "111111110101110101",  "111111110101110011",  "111111110101110000",  "111111110101101110",  "111111110101101011",  "111111110101101001",  "111111110101100110",  "111111110101100100",  "111111110101100001",  "111111110101011111",  "111111110101011101",  "111111110101011010",  "111111110101011000",  "111111110101010101",  "111111110101010011",  "111111110101010001",  "111111110101001110",  "111111110101001100",  "111111110101001001",  "111111110101000111",  "111111110101000101",  "111111110101000010",  "111111110101000000",  "111111110100111110",  "111111110100111011",  "111111110100111001",  "111111110100110111",  "111111110100110100",  "111111110100110010",  "111111110100110000",  "111111110100101110",  "111111110100101011",  "111111110100101001",  "111111110100100111",  "111111110100100101",  "111111110100100010",  "111111110100100000",  "111111110100011110",  "111111110100011100",  "111111110100011001",  "111111110100010111",  "111111110100010101",  "111111110100010011",  "111111110100010001",  "111111110100001110",  "111111110100001100",  "111111110100001010",  "111111110100001000",  "111111110100000110",  "111111110100000100",  "111111110100000010",  "111111110100000000",  "111111110011111101",  "111111110011111011",  "111111110011111001",  "111111110011110111",  "111111110011110101",  "111111110011110011",  "111111110011110001",  "111111110011101111",  "111111110011101101",  "111111110011101011",  "111111110011101001",  "111111110011100111",  "111111110011100101",  "111111110011100011",  "111111110011100001",  "111111110011011111",  "111111110011011101",  "111111110011011011",  "111111110011011001",  "111111110011010111",  "111111110011010101",  "111111110011010011",  "111111110011010001",  "111111110011001111",  "111111110011001101",  "111111110011001011",  "111111110011001010",  "111111110011001000",  "111111110011000110",  "111111110011000100",  "111111110011000010",  "111111110011000000",  "111111110010111110",  "111111110010111101",  "111111110010111011",  "111111110010111001",  "111111110010110111",  "111111110010110101",  "111111110010110100",  "111111110010110010",  "111111110010110000",  "111111110010101110",  "111111110010101100",  "111111110010101011",  "111111110010101001",  "111111110010100111",  "111111110010100110",  "111111110010100100",  "111111110010100010",  "111111110010100000",  "111111110010011111",  "111111110010011101",  "111111110010011011",  "111111110010011010",  "111111110010011000",  "111111110010010110",  "111111110010010101",  "111111110010010011",  "111111110010010010",  "111111110010010000",  "111111110010001110",  "111111110010001101",  "111111110010001011",  "111111110010001010",  "111111110010001000",  "111111110010000111",  "111111110010000101",  "111111110010000100",  "111111110010000010",  "111111110010000000",  "111111110001111111",  "111111110001111101",  "111111110001111100",  "111111110001111011",  "111111110001111001",  "111111110001111000",  "111111110001110110",  "111111110001110101",  "111111110001110011",  "111111110001110010",  "111111110001110000",  "111111110001101111",  "111111110001101110",  "111111110001101100",  "111111110001101011",  "111111110001101010",  "111111110001101000",  "111111110001100111",  "111111110001100101",  "111111110001100100",  "111111110001100011",  "111111110001100001",  "111111110001100000",  "111111110001011111",  "111111110001011110",  "111111110001011100",  "111111110001011011",  "111111110001011010",  "111111110001011001",  "111111110001010111",  "111111110001010110",  "111111110001010101",  "111111110001010100",  "111111110001010010",  "111111110001010001",  "111111110001010000",  "111111110001001111",  "111111110001001110",  "111111110001001101",  "111111110001001011",  "111111110001001010",  "111111110001001001",  "111111110001001000",  "111111110001000111",  "111111110001000110",  "111111110001000101",  "111111110001000100",  "111111110001000011",  "111111110001000010",  "111111110001000001",  "111111110001000000",  "111111110000111111",  "111111110000111101",  "111111110000111100",  "111111110000111011",  "111111110000111010",  "111111110000111001",  "111111110000111001",  "111111110000111000",  "111111110000110111",  "111111110000110110",  "111111110000110101",  "111111110000110100",  "111111110000110011",  "111111110000110010",  "111111110000110001",  "111111110000110000",  "111111110000101111",  "111111110000101110",  "111111110000101110",  "111111110000101101",  "111111110000101100",  "111111110000101011",  "111111110000101010",  "111111110000101001",  "111111110000101001",  "111111110000101000",  "111111110000100111",  "111111110000100110",  "111111110000100110",  "111111110000100101",  "111111110000100100",  "111111110000100011",  "111111110000100011",  "111111110000100010",  "111111110000100001",  "111111110000100000",  "111111110000100000",  "111111110000011111",  "111111110000011110",  "111111110000011110",  "111111110000011101",  "111111110000011101",  "111111110000011100",  "111111110000011011",  "111111110000011011",  "111111110000011010",  "111111110000011001",  "111111110000011001",  "111111110000011000",  "111111110000011000",  "111111110000010111",  "111111110000010111",  "111111110000010110",  "111111110000010110",  "111111110000010101",  "111111110000010101",  "111111110000010100",  "111111110000010100",  "111111110000010011",  "111111110000010011",  "111111110000010010",  "111111110000010010",  "111111110000010001",  "111111110000010001",  "111111110000010001",  "111111110000010000",  "111111110000010000",  "111111110000001111",  "111111110000001111",  "111111110000001111",  "111111110000001110",  "111111110000001110",  "111111110000001110",  "111111110000001101",  "111111110000001101",  "111111110000001101",  "111111110000001100",  "111111110000001100",  "111111110000001100",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001000",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001001",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001010",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001011",  "111111110000001100",  "111111110000001100",  "111111110000001100",  "111111110000001100",  "111111110000001101",  "111111110000001101",  "111111110000001101",  "111111110000001110",  "111111110000001110",  "111111110000001110",  "111111110000001111",  "111111110000001111",  "111111110000001111",  "111111110000010000",  "111111110000010000",  "111111110000010001",  "111111110000010001",  "111111110000010001",  "111111110000010010",  "111111110000010010",  "111111110000010011",  "111111110000010011",  "111111110000010100",  "111111110000010100",  "111111110000010101",  "111111110000010101",  "111111110000010110",  "111111110000010110",  "111111110000010111",  "111111110000010111",  "111111110000011000",  "111111110000011000",  "111111110000011001",  "111111110000011001",  "111111110000011010",  "111111110000011011",  "111111110000011011",  "111111110000011100",  "111111110000011100",  "111111110000011101",  "111111110000011110",  "111111110000011110",  "111111110000011111",  "111111110000100000",  "111111110000100000",  "111111110000100001",  "111111110000100010",  "111111110000100010",  "111111110000100011",  "111111110000100100",  "111111110000100100",  "111111110000100101",  "111111110000100110",  "111111110000100111",  "111111110000100111",  "111111110000101000",  "111111110000101001",  "111111110000101010",  "111111110000101011",  "111111110000101011",  "111111110000101100",  "111111110000101101",  "111111110000101110",  "111111110000101111",  "111111110000101111",  "111111110000110000",  "111111110000110001",  "111111110000110010",  "111111110000110011",  "111111110000110100",  "111111110000110101",  "111111110000110110",  "111111110000110111",  "111111110000111000",  "111111110000111000",  "111111110000111001",  "111111110000111010",  "111111110000111011",  "111111110000111100",  "111111110000111101",  "111111110000111110",  "111111110000111111",  "111111110001000000",  "111111110001000001",  "111111110001000010",  "111111110001000011",  "111111110001000100",  "111111110001000101",  "111111110001000111",  "111111110001001000",  "111111110001001001",  "111111110001001010",  "111111110001001011",  "111111110001001100",  "111111110001001101",  "111111110001001110",  "111111110001001111",  "111111110001010000",  "111111110001010010",  "111111110001010011",  "111111110001010100",  "111111110001010101",  "111111110001010110",  "111111110001010111",  "111111110001011001",  "111111110001011010",  "111111110001011011",  "111111110001011100",  "111111110001011101",  "111111110001011111",  "111111110001100000",  "111111110001100001",  "111111110001100010",  "111111110001100100",  "111111110001100101",  "111111110001100110",  "111111110001101000",  "111111110001101001",  "111111110001101010",  "111111110001101100",  "111111110001101101",  "111111110001101110",  "111111110001110000",  "111111110001110001",  "111111110001110010",  "111111110001110100",  "111111110001110101",  "111111110001110110",  "111111110001111000",  "111111110001111001",  "111111110001111011",  "111111110001111100",  "111111110001111101",  "111111110001111111",  "111111110010000000",  "111111110010000010",  "111111110010000011",  "111111110010000101",  "111111110010000110",  "111111110010001000",  "111111110010001001",  "111111110010001011",  "111111110010001100",  "111111110010001110",  "111111110010001111",  "111111110010010001",  "111111110010010010",  "111111110010010100",  "111111110010010101",  "111111110010010111",  "111111110010011000",  "111111110010011010",  "111111110010011100",  "111111110010011101",  "111111110010011111",  "111111110010100000",  "111111110010100010",  "111111110010100100",  "111111110010100101",  "111111110010100111",  "111111110010101000",  "111111110010101010",  "111111110010101100",  "111111110010101101",  "111111110010101111",  "111111110010110001",  "111111110010110010",  "111111110010110100",  "111111110010110110",  "111111110010111000",  "111111110010111001",  "111111110010111011",  "111111110010111101",  "111111110010111110",  "111111110011000000",  "111111110011000010",  "111111110011000100",  "111111110011000101",  "111111110011000111",  "111111110011001001",  "111111110011001011",  "111111110011001101",  "111111110011001110",  "111111110011010000",  "111111110011010010",  "111111110011010100",  "111111110011010110",  "111111110011011000",  "111111110011011001",  "111111110011011011",  "111111110011011101",  "111111110011011111",  "111111110011100001",  "111111110011100011",  "111111110011100101",  "111111110011100110",  "111111110011101000",  "111111110011101010",  "111111110011101100",  "111111110011101110",  "111111110011110000",  "111111110011110010",  "111111110011110100",  "111111110011110110",  "111111110011111000",  "111111110011111010",  "111111110011111100",  "111111110011111110",  "111111110100000000",  "111111110100000010",  "111111110100000100",  "111111110100000110",  "111111110100001000",  "111111110100001010",  "111111110100001100",  "111111110100001110",  "111111110100010000",  "111111110100010010",  "111111110100010100",  "111111110100010110",  "111111110100011000",  "111111110100011010",  "111111110100011100",  "111111110100011110",  "111111110100100000",  "111111110100100010",  "111111110100100100",  "111111110100100110",  "111111110100101000",  "111111110100101011",  "111111110100101101",  "111111110100101111",  "111111110100110001",  "111111110100110011",  "111111110100110101",  "111111110100110111",  "111111110100111001",  "111111110100111100",  "111111110100111110",  "111111110101000000",  "111111110101000010",  "111111110101000100",  "111111110101000110",  "111111110101001001",  "111111110101001011",  "111111110101001101",  "111111110101001111",  "111111110101010001",  "111111110101010100",  "111111110101010110",  "111111110101011000",  "111111110101011010",  "111111110101011101",  "111111110101011111",  "111111110101100001",  "111111110101100011",  "111111110101100110",  "111111110101101000",  "111111110101101010",  "111111110101101100",  "111111110101101111",  "111111110101110001",  "111111110101110011",  "111111110101110110",  "111111110101111000",  "111111110101111010",  "111111110101111101",  "111111110101111111",  "111111110110000001",  "111111110110000100",  "111111110110000110",  "111111110110001000",  "111111110110001011",  "111111110110001101",  "111111110110001111",  "111111110110010010",  "111111110110010100",  "111111110110010110",  "111111110110011001",  "111111110110011011",  "111111110110011110",  "111111110110100000",  "111111110110100010",  "111111110110100101",  "111111110110100111",  "111111110110101010",  "111111110110101100",  "111111110110101110",  "111111110110110001",  "111111110110110011",  "111111110110110110",  "111111110110111000",  "111111110110111011",  "111111110110111101",  "111111110110111111",  "111111110111000010",  "111111110111000100",  "111111110111000111",  "111111110111001001",  "111111110111001100",  "111111110111001110",  "111111110111010001",  "111111110111010011",  "111111110111010110",  "111111110111011000",  "111111110111011011",  "111111110111011101",  "111111110111100000",  "111111110111100010",  "111111110111100101",  "111111110111100111",  "111111110111101010",  "111111110111101100",  "111111110111101111",  "111111110111110001",  "111111110111110100",  "111111110111110110",  "111111110111111001",  "111111110111111100",  "111111110111111110",  "111111111000000001",  "111111111000000011",  "111111111000000110",  "111111111000001000",  "111111111000001011",  "111111111000001101",  "111111111000010000",  "111111111000010011",  "111111111000010101",  "111111111000011000",  "111111111000011010",  "111111111000011101",  "111111111000100000",  "111111111000100010",  "111111111000100101",  "111111111000100111",  "111111111000101010",  "111111111000101101",  "111111111000101111",  "111111111000110010",  "111111111000110101",  "111111111000110111",  "111111111000111010",  "111111111000111101",  "111111111000111111",  "111111111001000010",  "111111111001000100",  "111111111001000111",  "111111111001001010",  "111111111001001100",  "111111111001001111",  "111111111001010010",  "111111111001010100",  "111111111001010111",  "111111111001011010",  "111111111001011100",  "111111111001011111",  "111111111001100010",  "111111111001100101",  "111111111001100111",  "111111111001101010",  "111111111001101101",  "111111111001101111",  "111111111001110010",  "111111111001110101",  "111111111001110111",  "111111111001111010",  "111111111001111101",  "111111111010000000",  "111111111010000010",  "111111111010000101",  "111111111010001000",  "111111111010001010",  "111111111010001101",  "111111111010010000",  "111111111010010011",  "111111111010010101",  "111111111010011000",  "111111111010011011",  "111111111010011110",  "111111111010100000",  "111111111010100011",  "111111111010100110",  "111111111010101001",  "111111111010101011",  "111111111010101110",  "111111111010110001",  "111111111010110100",  "111111111010110110",  "111111111010111001",  "111111111010111100",  "111111111010111111",  "111111111011000001",  "111111111011000100",  "111111111011000111",  "111111111011001010",  "111111111011001100",  "111111111011001111",  "111111111011010010",  "111111111011010101",  "111111111011011000",  "111111111011011010",  "111111111011011101",  "111111111011100000",  "111111111011100011",  "111111111011100110",  "111111111011101000",  "111111111011101011",  "111111111011101110",  "111111111011110001",  "111111111011110011",  "111111111011110110",  "111111111011111001",  "111111111011111100",  "111111111011111111",  "111111111100000001",  "111111111100000100",  "111111111100000111",  "111111111100001010",  "111111111100001101",  "111111111100010000",  "111111111100010010",  "111111111100010101",  "111111111100011000",  "111111111100011011",  "111111111100011110",  "111111111100100000",  "111111111100100011",  "111111111100100110",  "111111111100101001",  "111111111100101100",  "111111111100101111",  "111111111100110001",  "111111111100110100",  "111111111100110111",  "111111111100111010",  "111111111100111101",  "111111111100111111",  "111111111101000010",  "111111111101000101",  "111111111101001000",  "111111111101001011",  "111111111101001110",  "111111111101010000",  "111111111101010011",  "111111111101010110",  "111111111101011001",  "111111111101011100",  "111111111101011111",  "111111111101100001",  "111111111101100100",  "111111111101100111",  "111111111101101010",  "111111111101101101",  "111111111101110000",  "111111111101110010",  "111111111101110101",  "111111111101111000",  "111111111101111011",  "111111111101111110",  "111111111110000001",  "111111111110000100",  "111111111110000110",  "111111111110001001",  "111111111110001100",  "111111111110001111",  "111111111110010010",  "111111111110010101",  "111111111110010111",  "111111111110011010",  "111111111110011101",  "111111111110100000",  "111111111110100011",  "111111111110100110",  "111111111110101000",  "111111111110101011",  "111111111110101110",  "111111111110110001",  "111111111110110100",  "111111111110110111",  "111111111110111001",  "111111111110111100",  "111111111110111111",  "111111111111000010",  "111111111111000101",  "111111111111001000",  "111111111111001010",  "111111111111001101",  "111111111111010000",  "111111111111010011",  "111111111111010110",  "111111111111011001",  "111111111111011011",  "111111111111011110",  "111111111111100001",  "111111111111100100",  "111111111111100111",  "111111111111101001",  "111111111111101100",  "111111111111101111",  "111111111111110010",  "111111111111110101",  "111111111111111000",  "111111111111111010",  "111111111111111101"),("000000000000000000",  "000000000000000011",  "000000000000000110",  "000000000000001000",  "000000000000001011",  "000000000000001110",  "000000000000010001",  "000000000000010100",  "000000000000010110",  "000000000000011001",  "000000000000011100",  "000000000000011111",  "000000000000100010",  "000000000000100100",  "000000000000100111",  "000000000000101010",  "000000000000101101",  "000000000000110000",  "000000000000110010",  "000000000000110101",  "000000000000111000",  "000000000000111011",  "000000000000111110",  "000000000001000000",  "000000000001000011",  "000000000001000110",  "000000000001001001",  "000000000001001011",  "000000000001001110",  "000000000001010001",  "000000000001010100",  "000000000001010111",  "000000000001011001",  "000000000001011100",  "000000000001011111",  "000000000001100010",  "000000000001100100",  "000000000001100111",  "000000000001101010",  "000000000001101101",  "000000000001101111",  "000000000001110010",  "000000000001110101",  "000000000001111000",  "000000000001111010",  "000000000001111101",  "000000000010000000",  "000000000010000011",  "000000000010000101",  "000000000010001000",  "000000000010001011",  "000000000010001101",  "000000000010010000",  "000000000010010011",  "000000000010010110",  "000000000010011000",  "000000000010011011",  "000000000010011110",  "000000000010100000",  "000000000010100011",  "000000000010100110",  "000000000010101001",  "000000000010101011",  "000000000010101110",  "000000000010110001",  "000000000010110011",  "000000000010110110",  "000000000010111001",  "000000000010111011",  "000000000010111110",  "000000000011000001",  "000000000011000011",  "000000000011000110",  "000000000011001001",  "000000000011001011",  "000000000011001110",  "000000000011010001",  "000000000011010011",  "000000000011010110",  "000000000011011001",  "000000000011011011",  "000000000011011110",  "000000000011100001",  "000000000011100011",  "000000000011100110",  "000000000011101000",  "000000000011101011",  "000000000011101110",  "000000000011110000",  "000000000011110011",  "000000000011110110",  "000000000011111000",  "000000000011111011",  "000000000011111101",  "000000000100000000",  "000000000100000011",  "000000000100000101",  "000000000100001000",  "000000000100001010",  "000000000100001101",  "000000000100010000",  "000000000100010010",  "000000000100010101",  "000000000100010111",  "000000000100011010",  "000000000100011100",  "000000000100011111",  "000000000100100001",  "000000000100100100",  "000000000100100111",  "000000000100101001",  "000000000100101100",  "000000000100101110",  "000000000100110001",  "000000000100110011",  "000000000100110110",  "000000000100111000",  "000000000100111011",  "000000000100111101",  "000000000101000000",  "000000000101000010",  "000000000101000101",  "000000000101000111",  "000000000101001010",  "000000000101001100",  "000000000101001111",  "000000000101010001",  "000000000101010100",  "000000000101010110",  "000000000101011001",  "000000000101011011",  "000000000101011110",  "000000000101100000",  "000000000101100010",  "000000000101100101",  "000000000101100111",  "000000000101101010",  "000000000101101100",  "000000000101101111",  "000000000101110001",  "000000000101110011",  "000000000101110110",  "000000000101111000",  "000000000101111011",  "000000000101111101",  "000000000101111111",  "000000000110000010",  "000000000110000100",  "000000000110000111",  "000000000110001001",  "000000000110001011",  "000000000110001110",  "000000000110010000",  "000000000110010010",  "000000000110010101",  "000000000110010111",  "000000000110011001",  "000000000110011100",  "000000000110011110",  "000000000110100000",  "000000000110100011",  "000000000110100101",  "000000000110100111",  "000000000110101010",  "000000000110101100",  "000000000110101110",  "000000000110110001",  "000000000110110011",  "000000000110110101",  "000000000110110111",  "000000000110111010",  "000000000110111100",  "000000000110111110",  "000000000111000000",  "000000000111000011",  "000000000111000101",  "000000000111000111",  "000000000111001001",  "000000000111001100",  "000000000111001110",  "000000000111010000",  "000000000111010010",  "000000000111010101",  "000000000111010111",  "000000000111011001",  "000000000111011011",  "000000000111011101",  "000000000111100000",  "000000000111100010",  "000000000111100100",  "000000000111100110",  "000000000111101000",  "000000000111101010",  "000000000111101101",  "000000000111101111",  "000000000111110001",  "000000000111110011",  "000000000111110101",  "000000000111110111",  "000000000111111001",  "000000000111111011",  "000000000111111110",  "000000001000000000",  "000000001000000010",  "000000001000000100",  "000000001000000110",  "000000001000001000",  "000000001000001010",  "000000001000001100",  "000000001000001110",  "000000001000010000",  "000000001000010010",  "000000001000010100",  "000000001000010110",  "000000001000011000",  "000000001000011010",  "000000001000011100",  "000000001000011110",  "000000001000100000",  "000000001000100010",  "000000001000100100",  "000000001000100110",  "000000001000101000",  "000000001000101010",  "000000001000101100",  "000000001000101110",  "000000001000110000",  "000000001000110010",  "000000001000110100",  "000000001000110110",  "000000001000111000",  "000000001000111010",  "000000001000111100",  "000000001000111110",  "000000001001000000",  "000000001001000010",  "000000001001000100",  "000000001001000101",  "000000001001000111",  "000000001001001001",  "000000001001001011",  "000000001001001101",  "000000001001001111",  "000000001001010001",  "000000001001010011",  "000000001001010100",  "000000001001010110",  "000000001001011000",  "000000001001011010",  "000000001001011100",  "000000001001011101",  "000000001001011111",  "000000001001100001",  "000000001001100011",  "000000001001100101",  "000000001001100110",  "000000001001101000",  "000000001001101010",  "000000001001101100",  "000000001001101101",  "000000001001101111",  "000000001001110001",  "000000001001110011",  "000000001001110100",  "000000001001110110",  "000000001001111000",  "000000001001111010",  "000000001001111011",  "000000001001111101",  "000000001001111111",  "000000001010000000",  "000000001010000010",  "000000001010000100",  "000000001010000101",  "000000001010000111",  "000000001010001001",  "000000001010001010",  "000000001010001100",  "000000001010001101",  "000000001010001111",  "000000001010010001",  "000000001010010010",  "000000001010010100",  "000000001010010101",  "000000001010010111",  "000000001010011001",  "000000001010011010",  "000000001010011100",  "000000001010011101",  "000000001010011111",  "000000001010100000",  "000000001010100010",  "000000001010100011",  "000000001010100101",  "000000001010100110",  "000000001010101000",  "000000001010101010",  "000000001010101011",  "000000001010101100",  "000000001010101110",  "000000001010101111",  "000000001010110001",  "000000001010110010",  "000000001010110100",  "000000001010110101",  "000000001010110111",  "000000001010111000",  "000000001010111010",  "000000001010111011",  "000000001010111100",  "000000001010111110",  "000000001010111111",  "000000001011000001",  "000000001011000010",  "000000001011000011",  "000000001011000101",  "000000001011000110",  "000000001011000111",  "000000001011001001",  "000000001011001010",  "000000001011001011",  "000000001011001101",  "000000001011001110",  "000000001011001111",  "000000001011010001",  "000000001011010010",  "000000001011010011",  "000000001011010100",  "000000001011010110",  "000000001011010111",  "000000001011011000",  "000000001011011001",  "000000001011011011",  "000000001011011100",  "000000001011011101",  "000000001011011110",  "000000001011100000",  "000000001011100001",  "000000001011100010",  "000000001011100011",  "000000001011100100",  "000000001011100101",  "000000001011100111",  "000000001011101000",  "000000001011101001",  "000000001011101010",  "000000001011101011",  "000000001011101100",  "000000001011101101",  "000000001011101111",  "000000001011110000",  "000000001011110001",  "000000001011110010",  "000000001011110011",  "000000001011110100",  "000000001011110101",  "000000001011110110",  "000000001011110111",  "000000001011111000",  "000000001011111001",  "000000001011111010",  "000000001011111011",  "000000001011111100",  "000000001011111101",  "000000001011111110",  "000000001011111111",  "000000001100000000",  "000000001100000001",  "000000001100000010",  "000000001100000011",  "000000001100000100",  "000000001100000101",  "000000001100000110",  "000000001100000111",  "000000001100001000",  "000000001100001001",  "000000001100001010",  "000000001100001011",  "000000001100001011",  "000000001100001100",  "000000001100001101",  "000000001100001110",  "000000001100001111",  "000000001100010000",  "000000001100010001",  "000000001100010001",  "000000001100010010",  "000000001100010011",  "000000001100010100",  "000000001100010101",  "000000001100010110",  "000000001100010110",  "000000001100010111",  "000000001100011000",  "000000001100011001",  "000000001100011001",  "000000001100011010",  "000000001100011011",  "000000001100011100",  "000000001100011100",  "000000001100011101",  "000000001100011110",  "000000001100011111",  "000000001100011111",  "000000001100100000",  "000000001100100001",  "000000001100100001",  "000000001100100010",  "000000001100100011",  "000000001100100011",  "000000001100100100",  "000000001100100100",  "000000001100100101",  "000000001100100110",  "000000001100100110",  "000000001100100111",  "000000001100101000",  "000000001100101000",  "000000001100101001",  "000000001100101001",  "000000001100101010",  "000000001100101010",  "000000001100101011",  "000000001100101011",  "000000001100101100",  "000000001100101100",  "000000001100101101",  "000000001100101110",  "000000001100101110",  "000000001100101111",  "000000001100101111",  "000000001100101111",  "000000001100110000",  "000000001100110000",  "000000001100110001",  "000000001100110001",  "000000001100110010",  "000000001100110010",  "000000001100110011",  "000000001100110011",  "000000001100110011",  "000000001100110100",  "000000001100110100",  "000000001100110101",  "000000001100110101",  "000000001100110101",  "000000001100110110",  "000000001100110110",  "000000001100110110",  "000000001100110111",  "000000001100110111",  "000000001100110111",  "000000001100111000",  "000000001100111000",  "000000001100111000",  "000000001100111000",  "000000001100111001",  "000000001100111001",  "000000001100111001",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111101",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111100",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111011",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111010",  "000000001100111001",  "000000001100111001",  "000000001100111001",  "000000001100111001",  "000000001100111000",  "000000001100111000",  "000000001100111000",  "000000001100110111",  "000000001100110111",  "000000001100110111",  "000000001100110110",  "000000001100110110",  "000000001100110110",  "000000001100110101",  "000000001100110101",  "000000001100110101",  "000000001100110100",  "000000001100110100",  "000000001100110100",  "000000001100110011",  "000000001100110011",  "000000001100110010",  "000000001100110010",  "000000001100110001",  "000000001100110001",  "000000001100110001",  "000000001100110000",  "000000001100110000",  "000000001100101111",  "000000001100101111",  "000000001100101110",  "000000001100101110",  "000000001100101101",  "000000001100101101",  "000000001100101100",  "000000001100101100",  "000000001100101011",  "000000001100101011",  "000000001100101010",  "000000001100101010",  "000000001100101001",  "000000001100101001",  "000000001100101000",  "000000001100100111",  "000000001100100111",  "000000001100100110",  "000000001100100110",  "000000001100100101",  "000000001100100100",  "000000001100100100",  "000000001100100011",  "000000001100100011",  "000000001100100010",  "000000001100100001",  "000000001100100001",  "000000001100100000",  "000000001100011111",  "000000001100011111",  "000000001100011110",  "000000001100011101",  "000000001100011101",  "000000001100011100",  "000000001100011011",  "000000001100011010",  "000000001100011010",  "000000001100011001",  "000000001100011000",  "000000001100010111",  "000000001100010111",  "000000001100010110",  "000000001100010101",  "000000001100010100",  "000000001100010100",  "000000001100010011",  "000000001100010010",  "000000001100010001",  "000000001100010000",  "000000001100010000",  "000000001100001111",  "000000001100001110",  "000000001100001101",  "000000001100001100",  "000000001100001011",  "000000001100001010",  "000000001100001010",  "000000001100001001",  "000000001100001000",  "000000001100000111",  "000000001100000110",  "000000001100000101",  "000000001100000100",  "000000001100000011",  "000000001100000010",  "000000001100000001",  "000000001100000001",  "000000001100000000",  "000000001011111111",  "000000001011111110",  "000000001011111101",  "000000001011111100",  "000000001011111011",  "000000001011111010",  "000000001011111001",  "000000001011111000",  "000000001011110111",  "000000001011110110",  "000000001011110101",  "000000001011110100",  "000000001011110011",  "000000001011110010",  "000000001011110001",  "000000001011101111",  "000000001011101110",  "000000001011101101",  "000000001011101100",  "000000001011101011",  "000000001011101010",  "000000001011101001",  "000000001011101000",  "000000001011100111",  "000000001011100110",  "000000001011100101",  "000000001011100011",  "000000001011100010",  "000000001011100001",  "000000001011100000",  "000000001011011111",  "000000001011011110",  "000000001011011101",  "000000001011011011",  "000000001011011010",  "000000001011011001",  "000000001011011000",  "000000001011010111",  "000000001011010101",  "000000001011010100",  "000000001011010011",  "000000001011010010",  "000000001011010001",  "000000001011001111",  "000000001011001110",  "000000001011001101",  "000000001011001100",  "000000001011001010",  "000000001011001001",  "000000001011001000",  "000000001011000110",  "000000001011000101",  "000000001011000100",  "000000001011000011",  "000000001011000001",  "000000001011000000",  "000000001010111111",  "000000001010111101",  "000000001010111100",  "000000001010111011",  "000000001010111001",  "000000001010111000",  "000000001010110111",  "000000001010110101",  "000000001010110100",  "000000001010110010",  "000000001010110001",  "000000001010110000",  "000000001010101110",  "000000001010101101",  "000000001010101100",  "000000001010101010",  "000000001010101001",  "000000001010100111",  "000000001010100110",  "000000001010100100",  "000000001010100011",  "000000001010100010",  "000000001010100000",  "000000001010011111",  "000000001010011101",  "000000001010011100",  "000000001010011010",  "000000001010011001",  "000000001010010111",  "000000001010010110",  "000000001010010100",  "000000001010010011",  "000000001010010001",  "000000001010010000",  "000000001010001110",  "000000001010001101",  "000000001010001011",  "000000001010001010",  "000000001010001000",  "000000001010000111",  "000000001010000101",  "000000001010000100",  "000000001010000010",  "000000001010000000",  "000000001001111111",  "000000001001111101",  "000000001001111100",  "000000001001111010",  "000000001001111000",  "000000001001110111",  "000000001001110101",  "000000001001110100",  "000000001001110010",  "000000001001110000",  "000000001001101111",  "000000001001101101",  "000000001001101100",  "000000001001101010",  "000000001001101000",  "000000001001100111",  "000000001001100101",  "000000001001100011",  "000000001001100010",  "000000001001100000",  "000000001001011110",  "000000001001011101",  "000000001001011011",  "000000001001011001",  "000000001001011000",  "000000001001010110",  "000000001001010100",  "000000001001010010",  "000000001001010001",  "000000001001001111",  "000000001001001101",  "000000001001001011",  "000000001001001010",  "000000001001001000",  "000000001001000110",  "000000001001000101",  "000000001001000011",  "000000001001000001",  "000000001000111111",  "000000001000111101",  "000000001000111100",  "000000001000111010",  "000000001000111000",  "000000001000110110",  "000000001000110101",  "000000001000110011",  "000000001000110001",  "000000001000101111",  "000000001000101101",  "000000001000101100",  "000000001000101010",  "000000001000101000",  "000000001000100110",  "000000001000100100",  "000000001000100010",  "000000001000100001",  "000000001000011111",  "000000001000011101",  "000000001000011011",  "000000001000011001",  "000000001000010111",  "000000001000010101",  "000000001000010100",  "000000001000010010",  "000000001000010000",  "000000001000001110",  "000000001000001100",  "000000001000001010",  "000000001000001000",  "000000001000000110",  "000000001000000100",  "000000001000000010",  "000000001000000001",  "000000000111111111",  "000000000111111101",  "000000000111111011",  "000000000111111001",  "000000000111110111",  "000000000111110101",  "000000000111110011",  "000000000111110001",  "000000000111101111",  "000000000111101101",  "000000000111101011",  "000000000111101001",  "000000000111100111",  "000000000111100101",  "000000000111100011",  "000000000111100001",  "000000000111011111",  "000000000111011101",  "000000000111011011",  "000000000111011001",  "000000000111010111",  "000000000111010101",  "000000000111010011",  "000000000111010001",  "000000000111001111",  "000000000111001101",  "000000000111001011",  "000000000111001001",  "000000000111000111",  "000000000111000101",  "000000000111000011",  "000000000111000001",  "000000000110111111",  "000000000110111101",  "000000000110111011",  "000000000110111001",  "000000000110110111",  "000000000110110101",  "000000000110110011",  "000000000110110001",  "000000000110101111",  "000000000110101101",  "000000000110101011",  "000000000110101001",  "000000000110100110",  "000000000110100100",  "000000000110100010",  "000000000110100000",  "000000000110011110",  "000000000110011100",  "000000000110011010",  "000000000110011000",  "000000000110010110",  "000000000110010100",  "000000000110010010",  "000000000110001111",  "000000000110001101",  "000000000110001011",  "000000000110001001",  "000000000110000111",  "000000000110000101",  "000000000110000011",  "000000000110000001",  "000000000101111110",  "000000000101111100",  "000000000101111010",  "000000000101111000",  "000000000101110110",  "000000000101110100",  "000000000101110010",  "000000000101101111",  "000000000101101101",  "000000000101101011",  "000000000101101001",  "000000000101100111",  "000000000101100101",  "000000000101100010",  "000000000101100000",  "000000000101011110",  "000000000101011100",  "000000000101011010",  "000000000101011000",  "000000000101010101",  "000000000101010011",  "000000000101010001",  "000000000101001111",  "000000000101001101",  "000000000101001010",  "000000000101001000",  "000000000101000110",  "000000000101000100",  "000000000101000010",  "000000000100111111",  "000000000100111101",  "000000000100111011",  "000000000100111001",  "000000000100110111",  "000000000100110100",  "000000000100110010",  "000000000100110000",  "000000000100101110",  "000000000100101100",  "000000000100101001",  "000000000100100111",  "000000000100100101",  "000000000100100011",  "000000000100100000",  "000000000100011110",  "000000000100011100",  "000000000100011010",  "000000000100010111",  "000000000100010101",  "000000000100010011",  "000000000100010001",  "000000000100001110",  "000000000100001100",  "000000000100001010",  "000000000100001000",  "000000000100000101",  "000000000100000011",  "000000000100000001",  "000000000011111111",  "000000000011111100",  "000000000011111010",  "000000000011111000",  "000000000011110110",  "000000000011110011",  "000000000011110001",  "000000000011101111",  "000000000011101101",  "000000000011101010",  "000000000011101000",  "000000000011100110",  "000000000011100100",  "000000000011100001",  "000000000011011111",  "000000000011011101",  "000000000011011010",  "000000000011011000",  "000000000011010110",  "000000000011010100",  "000000000011010001",  "000000000011001111",  "000000000011001101",  "000000000011001010",  "000000000011001000",  "000000000011000110",  "000000000011000100",  "000000000011000001",  "000000000010111111",  "000000000010111101",  "000000000010111010",  "000000000010111000",  "000000000010110110",  "000000000010110100",  "000000000010110001",  "000000000010101111",  "000000000010101101",  "000000000010101010",  "000000000010101000",  "000000000010100110",  "000000000010100011",  "000000000010100001",  "000000000010011111",  "000000000010011101",  "000000000010011010",  "000000000010011000",  "000000000010010110",  "000000000010010011",  "000000000010010001",  "000000000010001111",  "000000000010001100",  "000000000010001010",  "000000000010001000",  "000000000010000110",  "000000000010000011",  "000000000010000001",  "000000000001111111",  "000000000001111100",  "000000000001111010",  "000000000001111000",  "000000000001110101",  "000000000001110011",  "000000000001110001",  "000000000001101110",  "000000000001101100",  "000000000001101010",  "000000000001101000",  "000000000001100101",  "000000000001100011",  "000000000001100001",  "000000000001011110",  "000000000001011100",  "000000000001011010",  "000000000001010111",  "000000000001010101",  "000000000001010011",  "000000000001010000",  "000000000001001110",  "000000000001001100",  "000000000001001010",  "000000000001000111",  "000000000001000101",  "000000000001000011",  "000000000001000000",  "000000000000111110",  "000000000000111100",  "000000000000111001",  "000000000000110111",  "000000000000110101",  "000000000000110010",  "000000000000110000",  "000000000000101110",  "000000000000101100",  "000000000000101001",  "000000000000100111",  "000000000000100101",  "000000000000100010",  "000000000000100000",  "000000000000011110",  "000000000000011100",  "000000000000011001",  "000000000000010111",  "000000000000010101",  "000000000000010010",  "000000000000010000",  "000000000000001110",  "000000000000001011",  "000000000000001001",  "000000000000000111",  "000000000000000101",  "000000000000000010"),("000000000000000000",  "111111111111111110",  "111111111111111011",  "111111111111111001",  "111111111111110111",  "111111111111110101",  "111111111111110010",  "111111111111110000",  "111111111111101110",  "111111111111101011",  "111111111111101001",  "111111111111100111",  "111111111111100101",  "111111111111100010",  "111111111111100000",  "111111111111011110",  "111111111111011100",  "111111111111011001",  "111111111111010111",  "111111111111010101",  "111111111111010010",  "111111111111010000",  "111111111111001110",  "111111111111001100",  "111111111111001001",  "111111111111000111",  "111111111111000101",  "111111111111000011",  "111111111111000000",  "111111111110111110",  "111111111110111100",  "111111111110111010",  "111111111110110111",  "111111111110110101",  "111111111110110011",  "111111111110110001",  "111111111110101110",  "111111111110101100",  "111111111110101010",  "111111111110101000",  "111111111110100110",  "111111111110100011",  "111111111110100001",  "111111111110011111",  "111111111110011101",  "111111111110011010",  "111111111110011000",  "111111111110010110",  "111111111110010100",  "111111111110010010",  "111111111110001111",  "111111111110001101",  "111111111110001011",  "111111111110001001",  "111111111110000110",  "111111111110000100",  "111111111110000010",  "111111111110000000",  "111111111101111110",  "111111111101111011",  "111111111101111001",  "111111111101110111",  "111111111101110101",  "111111111101110011",  "111111111101110001",  "111111111101101110",  "111111111101101100",  "111111111101101010",  "111111111101101000",  "111111111101100110",  "111111111101100011",  "111111111101100001",  "111111111101011111",  "111111111101011101",  "111111111101011011",  "111111111101011001",  "111111111101010110",  "111111111101010100",  "111111111101010010",  "111111111101010000",  "111111111101001110",  "111111111101001100",  "111111111101001010",  "111111111101000111",  "111111111101000101",  "111111111101000011",  "111111111101000001",  "111111111100111111",  "111111111100111101",  "111111111100111011",  "111111111100111001",  "111111111100110110",  "111111111100110100",  "111111111100110010",  "111111111100110000",  "111111111100101110",  "111111111100101100",  "111111111100101010",  "111111111100101000",  "111111111100100110",  "111111111100100100",  "111111111100100001",  "111111111100011111",  "111111111100011101",  "111111111100011011",  "111111111100011001",  "111111111100010111",  "111111111100010101",  "111111111100010011",  "111111111100010001",  "111111111100001111",  "111111111100001101",  "111111111100001011",  "111111111100001001",  "111111111100000111",  "111111111100000101",  "111111111100000011",  "111111111100000000",  "111111111011111110",  "111111111011111100",  "111111111011111010",  "111111111011111000",  "111111111011110110",  "111111111011110100",  "111111111011110010",  "111111111011110000",  "111111111011101110",  "111111111011101100",  "111111111011101010",  "111111111011101000",  "111111111011100110",  "111111111011100100",  "111111111011100010",  "111111111011100000",  "111111111011011110",  "111111111011011100",  "111111111011011010",  "111111111011011000",  "111111111011010110",  "111111111011010100",  "111111111011010011",  "111111111011010001",  "111111111011001111",  "111111111011001101",  "111111111011001011",  "111111111011001001",  "111111111011000111",  "111111111011000101",  "111111111011000011",  "111111111011000001",  "111111111010111111",  "111111111010111101",  "111111111010111011",  "111111111010111001",  "111111111010111000",  "111111111010110110",  "111111111010110100",  "111111111010110010",  "111111111010110000",  "111111111010101110",  "111111111010101100",  "111111111010101010",  "111111111010101000",  "111111111010100111",  "111111111010100101",  "111111111010100011",  "111111111010100001",  "111111111010011111",  "111111111010011101",  "111111111010011011",  "111111111010011010",  "111111111010011000",  "111111111010010110",  "111111111010010100",  "111111111010010010",  "111111111010010000",  "111111111010001111",  "111111111010001101",  "111111111010001011",  "111111111010001001",  "111111111010000111",  "111111111010000110",  "111111111010000100",  "111111111010000010",  "111111111010000000",  "111111111001111110",  "111111111001111101",  "111111111001111011",  "111111111001111001",  "111111111001110111",  "111111111001110110",  "111111111001110100",  "111111111001110010",  "111111111001110000",  "111111111001101111",  "111111111001101101",  "111111111001101011",  "111111111001101001",  "111111111001101000",  "111111111001100110",  "111111111001100100",  "111111111001100011",  "111111111001100001",  "111111111001011111",  "111111111001011110",  "111111111001011100",  "111111111001011010",  "111111111001011001",  "111111111001010111",  "111111111001010101",  "111111111001010100",  "111111111001010010",  "111111111001010000",  "111111111001001111",  "111111111001001101",  "111111111001001011",  "111111111001001010",  "111111111001001000",  "111111111001000110",  "111111111001000101",  "111111111001000011",  "111111111001000010",  "111111111001000000",  "111111111000111110",  "111111111000111101",  "111111111000111011",  "111111111000111010",  "111111111000111000",  "111111111000110110",  "111111111000110101",  "111111111000110011",  "111111111000110010",  "111111111000110000",  "111111111000101111",  "111111111000101101",  "111111111000101100",  "111111111000101010",  "111111111000101000",  "111111111000100111",  "111111111000100101",  "111111111000100100",  "111111111000100010",  "111111111000100001",  "111111111000011111",  "111111111000011110",  "111111111000011100",  "111111111000011011",  "111111111000011001",  "111111111000011000",  "111111111000010110",  "111111111000010101",  "111111111000010100",  "111111111000010010",  "111111111000010001",  "111111111000001111",  "111111111000001110",  "111111111000001100",  "111111111000001011",  "111111111000001010",  "111111111000001000",  "111111111000000111",  "111111111000000101",  "111111111000000100",  "111111111000000010",  "111111111000000001",  "111111111000000000",  "111111110111111110",  "111111110111111101",  "111111110111111100",  "111111110111111010",  "111111110111111001",  "111111110111111000",  "111111110111110110",  "111111110111110101",  "111111110111110100",  "111111110111110010",  "111111110111110001",  "111111110111110000",  "111111110111101110",  "111111110111101101",  "111111110111101100",  "111111110111101010",  "111111110111101001",  "111111110111101000",  "111111110111100110",  "111111110111100101",  "111111110111100100",  "111111110111100011",  "111111110111100001",  "111111110111100000",  "111111110111011111",  "111111110111011110",  "111111110111011100",  "111111110111011011",  "111111110111011010",  "111111110111011001",  "111111110111011000",  "111111110111010110",  "111111110111010101",  "111111110111010100",  "111111110111010011",  "111111110111010010",  "111111110111010000",  "111111110111001111",  "111111110111001110",  "111111110111001101",  "111111110111001100",  "111111110111001011",  "111111110111001010",  "111111110111001000",  "111111110111000111",  "111111110111000110",  "111111110111000101",  "111111110111000100",  "111111110111000011",  "111111110111000010",  "111111110111000001",  "111111110111000000",  "111111110110111110",  "111111110110111101",  "111111110110111100",  "111111110110111011",  "111111110110111010",  "111111110110111001",  "111111110110111000",  "111111110110110111",  "111111110110110110",  "111111110110110101",  "111111110110110100",  "111111110110110011",  "111111110110110010",  "111111110110110001",  "111111110110110000",  "111111110110101111",  "111111110110101110",  "111111110110101101",  "111111110110101100",  "111111110110101011",  "111111110110101010",  "111111110110101001",  "111111110110101000",  "111111110110100111",  "111111110110100110",  "111111110110100101",  "111111110110100100",  "111111110110100100",  "111111110110100011",  "111111110110100010",  "111111110110100001",  "111111110110100000",  "111111110110011111",  "111111110110011110",  "111111110110011101",  "111111110110011100",  "111111110110011100",  "111111110110011011",  "111111110110011010",  "111111110110011001",  "111111110110011000",  "111111110110010111",  "111111110110010110",  "111111110110010110",  "111111110110010101",  "111111110110010100",  "111111110110010011",  "111111110110010010",  "111111110110010010",  "111111110110010001",  "111111110110010000",  "111111110110001111",  "111111110110001111",  "111111110110001110",  "111111110110001101",  "111111110110001100",  "111111110110001100",  "111111110110001011",  "111111110110001010",  "111111110110001001",  "111111110110001001",  "111111110110001000",  "111111110110000111",  "111111110110000111",  "111111110110000110",  "111111110110000101",  "111111110110000101",  "111111110110000100",  "111111110110000011",  "111111110110000011",  "111111110110000010",  "111111110110000001",  "111111110110000001",  "111111110110000000",  "111111110101111111",  "111111110101111111",  "111111110101111110",  "111111110101111101",  "111111110101111101",  "111111110101111100",  "111111110101111100",  "111111110101111011",  "111111110101111011",  "111111110101111010",  "111111110101111001",  "111111110101111001",  "111111110101111000",  "111111110101111000",  "111111110101110111",  "111111110101110111",  "111111110101110110",  "111111110101110110",  "111111110101110101",  "111111110101110101",  "111111110101110100",  "111111110101110100",  "111111110101110011",  "111111110101110011",  "111111110101110010",  "111111110101110010",  "111111110101110001",  "111111110101110001",  "111111110101110000",  "111111110101110000",  "111111110101101111",  "111111110101101111",  "111111110101101111",  "111111110101101110",  "111111110101101110",  "111111110101101101",  "111111110101101101",  "111111110101101101",  "111111110101101100",  "111111110101101100",  "111111110101101011",  "111111110101101011",  "111111110101101011",  "111111110101101010",  "111111110101101010",  "111111110101101010",  "111111110101101001",  "111111110101101001",  "111111110101101001",  "111111110101101000",  "111111110101101000",  "111111110101101000",  "111111110101101000",  "111111110101100111",  "111111110101100111",  "111111110101100111",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100001",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100010",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100011",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100100",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100101",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100110",  "111111110101100111",  "111111110101100111",  "111111110101100111",  "111111110101100111",  "111111110101101000",  "111111110101101000",  "111111110101101000",  "111111110101101001",  "111111110101101001",  "111111110101101001",  "111111110101101010",  "111111110101101010",  "111111110101101010",  "111111110101101011",  "111111110101101011",  "111111110101101011",  "111111110101101100",  "111111110101101100",  "111111110101101100",  "111111110101101101",  "111111110101101101",  "111111110101101110",  "111111110101101110",  "111111110101101110",  "111111110101101111",  "111111110101101111",  "111111110101110000",  "111111110101110000",  "111111110101110000",  "111111110101110001",  "111111110101110001",  "111111110101110010",  "111111110101110010",  "111111110101110011",  "111111110101110011",  "111111110101110100",  "111111110101110100",  "111111110101110101",  "111111110101110101",  "111111110101110110",  "111111110101110110",  "111111110101110111",  "111111110101110111",  "111111110101111000",  "111111110101111000",  "111111110101111001",  "111111110101111001",  "111111110101111010",  "111111110101111010",  "111111110101111011",  "111111110101111100",  "111111110101111100",  "111111110101111101",  "111111110101111101",  "111111110101111110",  "111111110101111110",  "111111110101111111",  "111111110110000000",  "111111110110000000",  "111111110110000001",  "111111110110000010",  "111111110110000010",  "111111110110000011",  "111111110110000011",  "111111110110000100",  "111111110110000101",  "111111110110000101",  "111111110110000110",  "111111110110000111",  "111111110110000111",  "111111110110001000",  "111111110110001001",  "111111110110001001",  "111111110110001010",  "111111110110001011",  "111111110110001100",  "111111110110001100",  "111111110110001101",  "111111110110001110",  "111111110110001110",  "111111110110001111",  "111111110110010000",  "111111110110010001",  "111111110110010001",  "111111110110010010",  "111111110110010011",  "111111110110010100",  "111111110110010101",  "111111110110010101",  "111111110110010110",  "111111110110010111",  "111111110110011000",  "111111110110011000",  "111111110110011001",  "111111110110011010",  "111111110110011011",  "111111110110011100",  "111111110110011101",  "111111110110011101",  "111111110110011110",  "111111110110011111",  "111111110110100000",  "111111110110100001",  "111111110110100010",  "111111110110100011",  "111111110110100011",  "111111110110100100",  "111111110110100101",  "111111110110100110",  "111111110110100111",  "111111110110101000",  "111111110110101001",  "111111110110101010",  "111111110110101011",  "111111110110101100",  "111111110110101100",  "111111110110101101",  "111111110110101110",  "111111110110101111",  "111111110110110000",  "111111110110110001",  "111111110110110010",  "111111110110110011",  "111111110110110100",  "111111110110110101",  "111111110110110110",  "111111110110110111",  "111111110110111000",  "111111110110111001",  "111111110110111010",  "111111110110111011",  "111111110110111100",  "111111110110111101",  "111111110110111110",  "111111110110111111",  "111111110111000000",  "111111110111000001",  "111111110111000010",  "111111110111000011",  "111111110111000100",  "111111110111000101",  "111111110111000110",  "111111110111000111",  "111111110111001001",  "111111110111001010",  "111111110111001011",  "111111110111001100",  "111111110111001101",  "111111110111001110",  "111111110111001111",  "111111110111010000",  "111111110111010001",  "111111110111010010",  "111111110111010011",  "111111110111010101",  "111111110111010110",  "111111110111010111",  "111111110111011000",  "111111110111011001",  "111111110111011010",  "111111110111011011",  "111111110111011101",  "111111110111011110",  "111111110111011111",  "111111110111100000",  "111111110111100001",  "111111110111100010",  "111111110111100100",  "111111110111100101",  "111111110111100110",  "111111110111100111",  "111111110111101000",  "111111110111101010",  "111111110111101011",  "111111110111101100",  "111111110111101101",  "111111110111101111",  "111111110111110000",  "111111110111110001",  "111111110111110010",  "111111110111110011",  "111111110111110101",  "111111110111110110",  "111111110111110111",  "111111110111111000",  "111111110111111010",  "111111110111111011",  "111111110111111100",  "111111110111111110",  "111111110111111111",  "111111111000000000",  "111111111000000001",  "111111111000000011",  "111111111000000100",  "111111111000000101",  "111111111000000111",  "111111111000001000",  "111111111000001001",  "111111111000001011",  "111111111000001100",  "111111111000001101",  "111111111000001111",  "111111111000010000",  "111111111000010001",  "111111111000010011",  "111111111000010100",  "111111111000010101",  "111111111000010111",  "111111111000011000",  "111111111000011001",  "111111111000011011",  "111111111000011100",  "111111111000011110",  "111111111000011111",  "111111111000100000",  "111111111000100010",  "111111111000100011",  "111111111000100100",  "111111111000100110",  "111111111000100111",  "111111111000101001",  "111111111000101010",  "111111111000101100",  "111111111000101101",  "111111111000101110",  "111111111000110000",  "111111111000110001",  "111111111000110011",  "111111111000110100",  "111111111000110110",  "111111111000110111",  "111111111000111000",  "111111111000111010",  "111111111000111011",  "111111111000111101",  "111111111000111110",  "111111111001000000",  "111111111001000001",  "111111111001000011",  "111111111001000100",  "111111111001000110",  "111111111001000111",  "111111111001001001",  "111111111001001010",  "111111111001001100",  "111111111001001101",  "111111111001001111",  "111111111001010000",  "111111111001010010",  "111111111001010011",  "111111111001010101",  "111111111001010110",  "111111111001011000",  "111111111001011001",  "111111111001011011",  "111111111001011100",  "111111111001011110",  "111111111001011111",  "111111111001100001",  "111111111001100011",  "111111111001100100",  "111111111001100110",  "111111111001100111",  "111111111001101001",  "111111111001101010",  "111111111001101100",  "111111111001101101",  "111111111001101111",  "111111111001110001",  "111111111001110010",  "111111111001110100",  "111111111001110101",  "111111111001110111",  "111111111001111001",  "111111111001111010",  "111111111001111100",  "111111111001111101",  "111111111001111111",  "111111111010000001",  "111111111010000010",  "111111111010000100",  "111111111010000101",  "111111111010000111",  "111111111010001001",  "111111111010001010",  "111111111010001100",  "111111111010001110",  "111111111010001111",  "111111111010010001",  "111111111010010010",  "111111111010010100",  "111111111010010110",  "111111111010010111",  "111111111010011001",  "111111111010011011",  "111111111010011100",  "111111111010011110",  "111111111010100000",  "111111111010100001",  "111111111010100011",  "111111111010100101",  "111111111010100110",  "111111111010101000",  "111111111010101010",  "111111111010101011",  "111111111010101101",  "111111111010101111",  "111111111010110000",  "111111111010110010",  "111111111010110100",  "111111111010110101",  "111111111010110111",  "111111111010111001",  "111111111010111011",  "111111111010111100",  "111111111010111110",  "111111111011000000",  "111111111011000001",  "111111111011000011",  "111111111011000101",  "111111111011000111",  "111111111011001000",  "111111111011001010",  "111111111011001100",  "111111111011001101",  "111111111011001111",  "111111111011010001",  "111111111011010011",  "111111111011010100",  "111111111011010110",  "111111111011011000",  "111111111011011010",  "111111111011011011",  "111111111011011101",  "111111111011011111",  "111111111011100001",  "111111111011100010",  "111111111011100100",  "111111111011100110",  "111111111011101000",  "111111111011101001",  "111111111011101011",  "111111111011101101",  "111111111011101111",  "111111111011110000",  "111111111011110010",  "111111111011110100",  "111111111011110110",  "111111111011110111",  "111111111011111001",  "111111111011111011",  "111111111011111101",  "111111111011111111",  "111111111100000000",  "111111111100000010",  "111111111100000100",  "111111111100000110",  "111111111100000111",  "111111111100001001",  "111111111100001011",  "111111111100001101",  "111111111100001111",  "111111111100010000",  "111111111100010010",  "111111111100010100",  "111111111100010110",  "111111111100011000",  "111111111100011001",  "111111111100011011",  "111111111100011101",  "111111111100011111",  "111111111100100001",  "111111111100100010",  "111111111100100100",  "111111111100100110",  "111111111100101000",  "111111111100101010",  "111111111100101100",  "111111111100101101",  "111111111100101111",  "111111111100110001",  "111111111100110011",  "111111111100110101",  "111111111100110110",  "111111111100111000",  "111111111100111010",  "111111111100111100",  "111111111100111110",  "111111111101000000",  "111111111101000001",  "111111111101000011",  "111111111101000101",  "111111111101000111",  "111111111101001001",  "111111111101001011",  "111111111101001100",  "111111111101001110",  "111111111101010000",  "111111111101010010",  "111111111101010100",  "111111111101010110",  "111111111101010111",  "111111111101011001",  "111111111101011011",  "111111111101011101",  "111111111101011111",  "111111111101100001",  "111111111101100010",  "111111111101100100",  "111111111101100110",  "111111111101101000",  "111111111101101010",  "111111111101101100",  "111111111101101110",  "111111111101101111",  "111111111101110001",  "111111111101110011",  "111111111101110101",  "111111111101110111",  "111111111101111001",  "111111111101111011",  "111111111101111100",  "111111111101111110",  "111111111110000000",  "111111111110000010",  "111111111110000100",  "111111111110000110",  "111111111110000111",  "111111111110001001",  "111111111110001011",  "111111111110001101",  "111111111110001111",  "111111111110010001",  "111111111110010011",  "111111111110010100",  "111111111110010110",  "111111111110011000",  "111111111110011010",  "111111111110011100",  "111111111110011110",  "111111111110100000",  "111111111110100001",  "111111111110100011",  "111111111110100101",  "111111111110100111",  "111111111110101001",  "111111111110101011",  "111111111110101101",  "111111111110101110",  "111111111110110000",  "111111111110110010",  "111111111110110100",  "111111111110110110",  "111111111110111000",  "111111111110111010",  "111111111110111100",  "111111111110111101",  "111111111110111111",  "111111111111000001",  "111111111111000011",  "111111111111000101",  "111111111111000111",  "111111111111001001",  "111111111111001010",  "111111111111001100",  "111111111111001110",  "111111111111010000",  "111111111111010010",  "111111111111010100",  "111111111111010101",  "111111111111010111",  "111111111111011001",  "111111111111011011",  "111111111111011101",  "111111111111011111",  "111111111111100001",  "111111111111100010",  "111111111111100100",  "111111111111100110",  "111111111111101000",  "111111111111101010",  "111111111111101100",  "111111111111101110",  "111111111111101111",  "111111111111110001",  "111111111111110011",  "111111111111110101",  "111111111111110111",  "111111111111111001",  "111111111111111010",  "111111111111111100",  "111111111111111110"),("000000000000000000",  "000000000000000010",  "000000000000000100",  "000000000000000110",  "000000000000000111",  "000000000000001001",  "000000000000001011",  "000000000000001101",  "000000000000001111",  "000000000000010001",  "000000000000010010",  "000000000000010100",  "000000000000010110",  "000000000000011000",  "000000000000011010",  "000000000000011100",  "000000000000011101",  "000000000000011111",  "000000000000100001",  "000000000000100011",  "000000000000100101",  "000000000000100110",  "000000000000101000",  "000000000000101010",  "000000000000101100",  "000000000000101110",  "000000000000110000",  "000000000000110001",  "000000000000110011",  "000000000000110101",  "000000000000110111",  "000000000000111001",  "000000000000111010",  "000000000000111100",  "000000000000111110",  "000000000001000000",  "000000000001000010",  "000000000001000011",  "000000000001000101",  "000000000001000111",  "000000000001001001",  "000000000001001011",  "000000000001001100",  "000000000001001110",  "000000000001010000",  "000000000001010010",  "000000000001010100",  "000000000001010101",  "000000000001010111",  "000000000001011001",  "000000000001011011",  "000000000001011100",  "000000000001011110",  "000000000001100000",  "000000000001100010",  "000000000001100100",  "000000000001100101",  "000000000001100111",  "000000000001101001",  "000000000001101011",  "000000000001101100",  "000000000001101110",  "000000000001110000",  "000000000001110010",  "000000000001110011",  "000000000001110101",  "000000000001110111",  "000000000001111001",  "000000000001111010",  "000000000001111100",  "000000000001111110",  "000000000010000000",  "000000000010000001",  "000000000010000011",  "000000000010000101",  "000000000010000111",  "000000000010001000",  "000000000010001010",  "000000000010001100",  "000000000010001110",  "000000000010001111",  "000000000010010001",  "000000000010010011",  "000000000010010100",  "000000000010010110",  "000000000010011000",  "000000000010011010",  "000000000010011011",  "000000000010011101",  "000000000010011111",  "000000000010100000",  "000000000010100010",  "000000000010100100",  "000000000010100101",  "000000000010100111",  "000000000010101001",  "000000000010101011",  "000000000010101100",  "000000000010101110",  "000000000010110000",  "000000000010110001",  "000000000010110011",  "000000000010110101",  "000000000010110110",  "000000000010111000",  "000000000010111010",  "000000000010111011",  "000000000010111101",  "000000000010111111",  "000000000011000000",  "000000000011000010",  "000000000011000100",  "000000000011000101",  "000000000011000111",  "000000000011001000",  "000000000011001010",  "000000000011001100",  "000000000011001101",  "000000000011001111",  "000000000011010001",  "000000000011010010",  "000000000011010100",  "000000000011010110",  "000000000011010111",  "000000000011011001",  "000000000011011010",  "000000000011011100",  "000000000011011110",  "000000000011011111",  "000000000011100001",  "000000000011100010",  "000000000011100100",  "000000000011100110",  "000000000011100111",  "000000000011101001",  "000000000011101010",  "000000000011101100",  "000000000011101110",  "000000000011101111",  "000000000011110001",  "000000000011110010",  "000000000011110100",  "000000000011110101",  "000000000011110111",  "000000000011111001",  "000000000011111010",  "000000000011111100",  "000000000011111101",  "000000000011111111",  "000000000100000000",  "000000000100000010",  "000000000100000011",  "000000000100000101",  "000000000100000110",  "000000000100001000",  "000000000100001001",  "000000000100001011",  "000000000100001101",  "000000000100001110",  "000000000100010000",  "000000000100010001",  "000000000100010011",  "000000000100010100",  "000000000100010110",  "000000000100010111",  "000000000100011001",  "000000000100011010",  "000000000100011100",  "000000000100011101",  "000000000100011110",  "000000000100100000",  "000000000100100001",  "000000000100100011",  "000000000100100100",  "000000000100100110",  "000000000100100111",  "000000000100101001",  "000000000100101010",  "000000000100101100",  "000000000100101101",  "000000000100101111",  "000000000100110000",  "000000000100110001",  "000000000100110011",  "000000000100110100",  "000000000100110110",  "000000000100110111",  "000000000100111001",  "000000000100111010",  "000000000100111011",  "000000000100111101",  "000000000100111110",  "000000000101000000",  "000000000101000001",  "000000000101000010",  "000000000101000100",  "000000000101000101",  "000000000101000110",  "000000000101001000",  "000000000101001001",  "000000000101001011",  "000000000101001100",  "000000000101001101",  "000000000101001111",  "000000000101010000",  "000000000101010001",  "000000000101010011",  "000000000101010100",  "000000000101010101",  "000000000101010111",  "000000000101011000",  "000000000101011001",  "000000000101011011",  "000000000101011100",  "000000000101011101",  "000000000101011111",  "000000000101100000",  "000000000101100001",  "000000000101100011",  "000000000101100100",  "000000000101100101",  "000000000101100110",  "000000000101101000",  "000000000101101001",  "000000000101101010",  "000000000101101100",  "000000000101101101",  "000000000101101110",  "000000000101101111",  "000000000101110001",  "000000000101110010",  "000000000101110011",  "000000000101110100",  "000000000101110110",  "000000000101110111",  "000000000101111000",  "000000000101111001",  "000000000101111011",  "000000000101111100",  "000000000101111101",  "000000000101111110",  "000000000101111111",  "000000000110000001",  "000000000110000010",  "000000000110000011",  "000000000110000100",  "000000000110000101",  "000000000110000111",  "000000000110001000",  "000000000110001001",  "000000000110001010",  "000000000110001011",  "000000000110001100",  "000000000110001110",  "000000000110001111",  "000000000110010000",  "000000000110010001",  "000000000110010010",  "000000000110010011",  "000000000110010100",  "000000000110010110",  "000000000110010111",  "000000000110011000",  "000000000110011001",  "000000000110011010",  "000000000110011011",  "000000000110011100",  "000000000110011101",  "000000000110011110",  "000000000110100000",  "000000000110100001",  "000000000110100010",  "000000000110100011",  "000000000110100100",  "000000000110100101",  "000000000110100110",  "000000000110100111",  "000000000110101000",  "000000000110101001",  "000000000110101010",  "000000000110101011",  "000000000110101100",  "000000000110101101",  "000000000110101110",  "000000000110101111",  "000000000110110000",  "000000000110110001",  "000000000110110010",  "000000000110110011",  "000000000110110100",  "000000000110110101",  "000000000110110110",  "000000000110110111",  "000000000110111000",  "000000000110111001",  "000000000110111010",  "000000000110111011",  "000000000110111100",  "000000000110111101",  "000000000110111110",  "000000000110111111",  "000000000111000000",  "000000000111000001",  "000000000111000010",  "000000000111000011",  "000000000111000100",  "000000000111000101",  "000000000111000110",  "000000000111000110",  "000000000111000111",  "000000000111001000",  "000000000111001001",  "000000000111001010",  "000000000111001011",  "000000000111001100",  "000000000111001101",  "000000000111001110",  "000000000111001110",  "000000000111001111",  "000000000111010000",  "000000000111010001",  "000000000111010010",  "000000000111010011",  "000000000111010011",  "000000000111010100",  "000000000111010101",  "000000000111010110",  "000000000111010111",  "000000000111011000",  "000000000111011000",  "000000000111011001",  "000000000111011010",  "000000000111011011",  "000000000111011100",  "000000000111011100",  "000000000111011101",  "000000000111011110",  "000000000111011111",  "000000000111011111",  "000000000111100000",  "000000000111100001",  "000000000111100010",  "000000000111100011",  "000000000111100011",  "000000000111100100",  "000000000111100101",  "000000000111100101",  "000000000111100110",  "000000000111100111",  "000000000111101000",  "000000000111101000",  "000000000111101001",  "000000000111101010",  "000000000111101010",  "000000000111101011",  "000000000111101100",  "000000000111101100",  "000000000111101101",  "000000000111101110",  "000000000111101110",  "000000000111101111",  "000000000111110000",  "000000000111110000",  "000000000111110001",  "000000000111110010",  "000000000111110010",  "000000000111110011",  "000000000111110100",  "000000000111110100",  "000000000111110101",  "000000000111110101",  "000000000111110110",  "000000000111110111",  "000000000111110111",  "000000000111111000",  "000000000111111000",  "000000000111111001",  "000000000111111010",  "000000000111111010",  "000000000111111011",  "000000000111111011",  "000000000111111100",  "000000000111111100",  "000000000111111101",  "000000000111111101",  "000000000111111110",  "000000000111111110",  "000000000111111111",  "000000000111111111",  "000000001000000000",  "000000001000000000",  "000000001000000001",  "000000001000000001",  "000000001000000010",  "000000001000000010",  "000000001000000011",  "000000001000000011",  "000000001000000100",  "000000001000000100",  "000000001000000101",  "000000001000000101",  "000000001000000110",  "000000001000000110",  "000000001000000111",  "000000001000000111",  "000000001000000111",  "000000001000001000",  "000000001000001000",  "000000001000001001",  "000000001000001001",  "000000001000001010",  "000000001000001010",  "000000001000001010",  "000000001000001011",  "000000001000001011",  "000000001000001011",  "000000001000001100",  "000000001000001100",  "000000001000001101",  "000000001000001101",  "000000001000001101",  "000000001000001110",  "000000001000001110",  "000000001000001110",  "000000001000001111",  "000000001000001111",  "000000001000001111",  "000000001000010000",  "000000001000010000",  "000000001000010000",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010010",  "000000001000010010",  "000000001000010010",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011001",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000011000",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010111",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010110",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010101",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010100",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010011",  "000000001000010010",  "000000001000010010",  "000000001000010010",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010001",  "000000001000010000",  "000000001000010000",  "000000001000010000",  "000000001000001111",  "000000001000001111",  "000000001000001111",  "000000001000001110",  "000000001000001110",  "000000001000001110",  "000000001000001101",  "000000001000001101",  "000000001000001101",  "000000001000001100",  "000000001000001100",  "000000001000001100",  "000000001000001011",  "000000001000001011",  "000000001000001011",  "000000001000001010",  "000000001000001010",  "000000001000001001",  "000000001000001001",  "000000001000001001",  "000000001000001000",  "000000001000001000",  "000000001000000111",  "000000001000000111",  "000000001000000111",  "000000001000000110",  "000000001000000110",  "000000001000000101",  "000000001000000101",  "000000001000000100",  "000000001000000100",  "000000001000000011",  "000000001000000011",  "000000001000000010",  "000000001000000010",  "000000001000000010",  "000000001000000001",  "000000001000000001",  "000000001000000000",  "000000001000000000",  "000000000111111111",  "000000000111111111",  "000000000111111110",  "000000000111111110",  "000000000111111101",  "000000000111111101",  "000000000111111100",  "000000000111111011",  "000000000111111011",  "000000000111111010",  "000000000111111010",  "000000000111111001",  "000000000111111001",  "000000000111111000",  "000000000111111000",  "000000000111110111",  "000000000111110110",  "000000000111110110",  "000000000111110101",  "000000000111110101",  "000000000111110100",  "000000000111110100",  "000000000111110011",  "000000000111110010",  "000000000111110010",  "000000000111110001",  "000000000111110000",  "000000000111110000",  "000000000111101111",  "000000000111101111",  "000000000111101110",  "000000000111101101",  "000000000111101101",  "000000000111101100",  "000000000111101011",  "000000000111101011",  "000000000111101010",  "000000000111101001",  "000000000111101001",  "000000000111101000",  "000000000111100111",  "000000000111100111",  "000000000111100110",  "000000000111100101",  "000000000111100101",  "000000000111100100",  "000000000111100011",  "000000000111100011",  "000000000111100010",  "000000000111100001",  "000000000111100000",  "000000000111100000",  "000000000111011111",  "000000000111011110",  "000000000111011101",  "000000000111011101",  "000000000111011100",  "000000000111011011",  "000000000111011010",  "000000000111011010",  "000000000111011001",  "000000000111011000",  "000000000111010111",  "000000000111010111",  "000000000111010110",  "000000000111010101",  "000000000111010100",  "000000000111010011",  "000000000111010011",  "000000000111010010",  "000000000111010001",  "000000000111010000",  "000000000111001111",  "000000000111001111",  "000000000111001110",  "000000000111001101",  "000000000111001100",  "000000000111001011",  "000000000111001010",  "000000000111001010",  "000000000111001001",  "000000000111001000",  "000000000111000111",  "000000000111000110",  "000000000111000101",  "000000000111000101",  "000000000111000100",  "000000000111000011",  "000000000111000010",  "000000000111000001",  "000000000111000000",  "000000000110111111",  "000000000110111110",  "000000000110111101",  "000000000110111101",  "000000000110111100",  "000000000110111011",  "000000000110111010",  "000000000110111001",  "000000000110111000",  "000000000110110111",  "000000000110110110",  "000000000110110101",  "000000000110110100",  "000000000110110011",  "000000000110110010",  "000000000110110001",  "000000000110110001",  "000000000110110000",  "000000000110101111",  "000000000110101110",  "000000000110101101",  "000000000110101100",  "000000000110101011",  "000000000110101010",  "000000000110101001",  "000000000110101000",  "000000000110100111",  "000000000110100110",  "000000000110100101",  "000000000110100100",  "000000000110100011",  "000000000110100010",  "000000000110100001",  "000000000110100000",  "000000000110011111",  "000000000110011110",  "000000000110011101",  "000000000110011100",  "000000000110011011",  "000000000110011010",  "000000000110011001",  "000000000110011000",  "000000000110010111",  "000000000110010110",  "000000000110010101",  "000000000110010011",  "000000000110010010",  "000000000110010001",  "000000000110010000",  "000000000110001111",  "000000000110001110",  "000000000110001101",  "000000000110001100",  "000000000110001011",  "000000000110001010",  "000000000110001001",  "000000000110001000",  "000000000110000111",  "000000000110000110",  "000000000110000100",  "000000000110000011",  "000000000110000010",  "000000000110000001",  "000000000110000000",  "000000000101111111",  "000000000101111110",  "000000000101111101",  "000000000101111100",  "000000000101111010",  "000000000101111001",  "000000000101111000",  "000000000101110111",  "000000000101110110",  "000000000101110101",  "000000000101110100",  "000000000101110011",  "000000000101110001",  "000000000101110000",  "000000000101101111",  "000000000101101110",  "000000000101101101",  "000000000101101100",  "000000000101101010",  "000000000101101001",  "000000000101101000",  "000000000101100111",  "000000000101100110",  "000000000101100101",  "000000000101100011",  "000000000101100010",  "000000000101100001",  "000000000101100000",  "000000000101011111",  "000000000101011101",  "000000000101011100",  "000000000101011011",  "000000000101011010",  "000000000101011001",  "000000000101010111",  "000000000101010110",  "000000000101010101",  "000000000101010100",  "000000000101010011",  "000000000101010001",  "000000000101010000",  "000000000101001111",  "000000000101001110",  "000000000101001100",  "000000000101001011",  "000000000101001010",  "000000000101001001",  "000000000101000111",  "000000000101000110",  "000000000101000101",  "000000000101000100",  "000000000101000010",  "000000000101000001",  "000000000101000000",  "000000000100111111",  "000000000100111101",  "000000000100111100",  "000000000100111011",  "000000000100111010",  "000000000100111000",  "000000000100110111",  "000000000100110110",  "000000000100110100",  "000000000100110011",  "000000000100110010",  "000000000100110001",  "000000000100101111",  "000000000100101110",  "000000000100101101",  "000000000100101011",  "000000000100101010",  "000000000100101001",  "000000000100100111",  "000000000100100110",  "000000000100100101",  "000000000100100100",  "000000000100100010",  "000000000100100001",  "000000000100100000",  "000000000100011110",  "000000000100011101",  "000000000100011100",  "000000000100011010",  "000000000100011001",  "000000000100011000",  "000000000100010110",  "000000000100010101",  "000000000100010100",  "000000000100010010",  "000000000100010001",  "000000000100010000",  "000000000100001110",  "000000000100001101",  "000000000100001100",  "000000000100001010",  "000000000100001001",  "000000000100001000",  "000000000100000110",  "000000000100000101",  "000000000100000011",  "000000000100000010",  "000000000100000001",  "000000000011111111",  "000000000011111110",  "000000000011111101",  "000000000011111011",  "000000000011111010",  "000000000011111001",  "000000000011110111",  "000000000011110110",  "000000000011110100",  "000000000011110011",  "000000000011110010",  "000000000011110000",  "000000000011101111",  "000000000011101110",  "000000000011101100",  "000000000011101011",  "000000000011101001",  "000000000011101000",  "000000000011100111",  "000000000011100101",  "000000000011100100",  "000000000011100010",  "000000000011100001",  "000000000011100000",  "000000000011011110",  "000000000011011101",  "000000000011011011",  "000000000011011010",  "000000000011011001",  "000000000011010111",  "000000000011010110",  "000000000011010100",  "000000000011010011",  "000000000011010001",  "000000000011010000",  "000000000011001111",  "000000000011001101",  "000000000011001100",  "000000000011001010",  "000000000011001001",  "000000000011000111",  "000000000011000110",  "000000000011000101",  "000000000011000011",  "000000000011000010",  "000000000011000000",  "000000000010111111",  "000000000010111101",  "000000000010111100",  "000000000010111011",  "000000000010111001",  "000000000010111000",  "000000000010110110",  "000000000010110101",  "000000000010110011",  "000000000010110010",  "000000000010110001",  "000000000010101111",  "000000000010101110",  "000000000010101100",  "000000000010101011",  "000000000010101001",  "000000000010101000",  "000000000010100110",  "000000000010100101",  "000000000010100011",  "000000000010100010",  "000000000010100001",  "000000000010011111",  "000000000010011110",  "000000000010011100",  "000000000010011011",  "000000000010011001",  "000000000010011000",  "000000000010010110",  "000000000010010101",  "000000000010010011",  "000000000010010010",  "000000000010010001",  "000000000010001111",  "000000000010001110",  "000000000010001100",  "000000000010001011",  "000000000010001001",  "000000000010001000",  "000000000010000110",  "000000000010000101",  "000000000010000011",  "000000000010000010",  "000000000010000000",  "000000000001111111",  "000000000001111101",  "000000000001111100",  "000000000001111011",  "000000000001111001",  "000000000001111000",  "000000000001110110",  "000000000001110101",  "000000000001110011",  "000000000001110010",  "000000000001110000",  "000000000001101111",  "000000000001101101",  "000000000001101100",  "000000000001101010",  "000000000001101001",  "000000000001100111",  "000000000001100110",  "000000000001100100",  "000000000001100011",  "000000000001100001",  "000000000001100000",  "000000000001011110",  "000000000001011101",  "000000000001011100",  "000000000001011010",  "000000000001011001",  "000000000001010111",  "000000000001010110",  "000000000001010100",  "000000000001010011",  "000000000001010001",  "000000000001010000",  "000000000001001110",  "000000000001001101",  "000000000001001011",  "000000000001001010",  "000000000001001000",  "000000000001000111",  "000000000001000101",  "000000000001000100",  "000000000001000010",  "000000000001000001",  "000000000000111111",  "000000000000111110",  "000000000000111100",  "000000000000111011",  "000000000000111001",  "000000000000111000",  "000000000000110111",  "000000000000110101",  "000000000000110100",  "000000000000110010",  "000000000000110001",  "000000000000101111",  "000000000000101110",  "000000000000101100",  "000000000000101011",  "000000000000101001",  "000000000000101000",  "000000000000100110",  "000000000000100101",  "000000000000100011",  "000000000000100010",  "000000000000100000",  "000000000000011111",  "000000000000011101",  "000000000000011100",  "000000000000011010",  "000000000000011001",  "000000000000011000",  "000000000000010110",  "000000000000010101",  "000000000000010011",  "000000000000010010",  "000000000000010000",  "000000000000001111",  "000000000000001101",  "000000000000001100",  "000000000000001010",  "000000000000001001",  "000000000000000111",  "000000000000000110",  "000000000000000100",  "000000000000000011",  "000000000000000001"),("000000000000000000",  "111111111111111111",  "111111111111111101",  "111111111111111100",  "111111111111111010",  "111111111111111001",  "111111111111110111",  "111111111111110110",  "111111111111110100",  "111111111111110011",  "111111111111110001",  "111111111111110000",  "111111111111101110",  "111111111111101101",  "111111111111101100",  "111111111111101010",  "111111111111101001",  "111111111111100111",  "111111111111100110",  "111111111111100100",  "111111111111100011",  "111111111111100001",  "111111111111100000",  "111111111111011111",  "111111111111011101",  "111111111111011100",  "111111111111011010",  "111111111111011001",  "111111111111010111",  "111111111111010110",  "111111111111010100",  "111111111111010011",  "111111111111010010",  "111111111111010000",  "111111111111001111",  "111111111111001101",  "111111111111001100",  "111111111111001010",  "111111111111001001",  "111111111111001000",  "111111111111000110",  "111111111111000101",  "111111111111000011",  "111111111111000010",  "111111111111000000",  "111111111110111111",  "111111111110111110",  "111111111110111100",  "111111111110111011",  "111111111110111001",  "111111111110111000",  "111111111110110111",  "111111111110110101",  "111111111110110100",  "111111111110110010",  "111111111110110001",  "111111111110101111",  "111111111110101110",  "111111111110101101",  "111111111110101011",  "111111111110101010",  "111111111110101000",  "111111111110100111",  "111111111110100110",  "111111111110100100",  "111111111110100011",  "111111111110100001",  "111111111110100000",  "111111111110011111",  "111111111110011101",  "111111111110011100",  "111111111110011011",  "111111111110011001",  "111111111110011000",  "111111111110010110",  "111111111110010101",  "111111111110010100",  "111111111110010010",  "111111111110010001",  "111111111110010000",  "111111111110001110",  "111111111110001101",  "111111111110001011",  "111111111110001010",  "111111111110001001",  "111111111110000111",  "111111111110000110",  "111111111110000101",  "111111111110000011",  "111111111110000010",  "111111111110000001",  "111111111101111111",  "111111111101111110",  "111111111101111101",  "111111111101111011",  "111111111101111010",  "111111111101111001",  "111111111101110111",  "111111111101110110",  "111111111101110100",  "111111111101110011",  "111111111101110010",  "111111111101110001",  "111111111101101111",  "111111111101101110",  "111111111101101101",  "111111111101101011",  "111111111101101010",  "111111111101101001",  "111111111101100111",  "111111111101100110",  "111111111101100101",  "111111111101100011",  "111111111101100010",  "111111111101100001",  "111111111101011111",  "111111111101011110",  "111111111101011101",  "111111111101011100",  "111111111101011010",  "111111111101011001",  "111111111101011000",  "111111111101010110",  "111111111101010101",  "111111111101010100",  "111111111101010011",  "111111111101010001",  "111111111101010000",  "111111111101001111",  "111111111101001101",  "111111111101001100",  "111111111101001011",  "111111111101001010",  "111111111101001000",  "111111111101000111",  "111111111101000110",  "111111111101000101",  "111111111101000011",  "111111111101000010",  "111111111101000001",  "111111111101000000",  "111111111100111110",  "111111111100111101",  "111111111100111100",  "111111111100111011",  "111111111100111001",  "111111111100111000",  "111111111100110111",  "111111111100110110",  "111111111100110100",  "111111111100110011",  "111111111100110010",  "111111111100110001",  "111111111100110000",  "111111111100101110",  "111111111100101101",  "111111111100101100",  "111111111100101011",  "111111111100101010",  "111111111100101000",  "111111111100100111",  "111111111100100110",  "111111111100100101",  "111111111100100100",  "111111111100100010",  "111111111100100001",  "111111111100100000",  "111111111100011111",  "111111111100011110",  "111111111100011101",  "111111111100011011",  "111111111100011010",  "111111111100011001",  "111111111100011000",  "111111111100010111",  "111111111100010110",  "111111111100010100",  "111111111100010011",  "111111111100010010",  "111111111100010001",  "111111111100010000",  "111111111100001111",  "111111111100001110",  "111111111100001100",  "111111111100001011",  "111111111100001010",  "111111111100001001",  "111111111100001000",  "111111111100000111",  "111111111100000110",  "111111111100000101",  "111111111100000011",  "111111111100000010",  "111111111100000001",  "111111111100000000",  "111111111011111111",  "111111111011111110",  "111111111011111101",  "111111111011111100",  "111111111011111011",  "111111111011111010",  "111111111011111001",  "111111111011110111",  "111111111011110110",  "111111111011110101",  "111111111011110100",  "111111111011110011",  "111111111011110010",  "111111111011110001",  "111111111011110000",  "111111111011101111",  "111111111011101110",  "111111111011101101",  "111111111011101100",  "111111111011101011",  "111111111011101010",  "111111111011101001",  "111111111011101000",  "111111111011100111",  "111111111011100110",  "111111111011100101",  "111111111011100100",  "111111111011100011",  "111111111011100010",  "111111111011100001",  "111111111011100000",  "111111111011011111",  "111111111011011110",  "111111111011011101",  "111111111011011100",  "111111111011011011",  "111111111011011010",  "111111111011011001",  "111111111011011000",  "111111111011010111",  "111111111011010110",  "111111111011010101",  "111111111011010100",  "111111111011010011",  "111111111011010010",  "111111111011010001",  "111111111011010000",  "111111111011001111",  "111111111011001110",  "111111111011001101",  "111111111011001100",  "111111111011001011",  "111111111011001010",  "111111111011001001",  "111111111011001000",  "111111111011000111",  "111111111011000111",  "111111111011000110",  "111111111011000101",  "111111111011000100",  "111111111011000011",  "111111111011000010",  "111111111011000001",  "111111111011000000",  "111111111010111111",  "111111111010111110",  "111111111010111101",  "111111111010111101",  "111111111010111100",  "111111111010111011",  "111111111010111010",  "111111111010111001",  "111111111010111000",  "111111111010110111",  "111111111010110111",  "111111111010110110",  "111111111010110101",  "111111111010110100",  "111111111010110011",  "111111111010110010",  "111111111010110001",  "111111111010110001",  "111111111010110000",  "111111111010101111",  "111111111010101110",  "111111111010101101",  "111111111010101101",  "111111111010101100",  "111111111010101011",  "111111111010101010",  "111111111010101001",  "111111111010101000",  "111111111010101000",  "111111111010100111",  "111111111010100110",  "111111111010100101",  "111111111010100101",  "111111111010100100",  "111111111010100011",  "111111111010100010",  "111111111010100001",  "111111111010100001",  "111111111010100000",  "111111111010011111",  "111111111010011110",  "111111111010011110",  "111111111010011101",  "111111111010011100",  "111111111010011011",  "111111111010011011",  "111111111010011010",  "111111111010011001",  "111111111010011001",  "111111111010011000",  "111111111010010111",  "111111111010010110",  "111111111010010110",  "111111111010010101",  "111111111010010100",  "111111111010010100",  "111111111010010011",  "111111111010010010",  "111111111010010010",  "111111111010010001",  "111111111010010000",  "111111111010010000",  "111111111010001111",  "111111111010001110",  "111111111010001110",  "111111111010001101",  "111111111010001100",  "111111111010001100",  "111111111010001011",  "111111111010001010",  "111111111010001010",  "111111111010001001",  "111111111010001000",  "111111111010001000",  "111111111010000111",  "111111111010000111",  "111111111010000110",  "111111111010000101",  "111111111010000101",  "111111111010000100",  "111111111010000100",  "111111111010000011",  "111111111010000010",  "111111111010000010",  "111111111010000001",  "111111111010000001",  "111111111010000000",  "111111111001111111",  "111111111001111111",  "111111111001111110",  "111111111001111110",  "111111111001111101",  "111111111001111101",  "111111111001111100",  "111111111001111100",  "111111111001111011",  "111111111001111011",  "111111111001111010",  "111111111001111001",  "111111111001111001",  "111111111001111000",  "111111111001111000",  "111111111001110111",  "111111111001110111",  "111111111001110110",  "111111111001110110",  "111111111001110101",  "111111111001110101",  "111111111001110100",  "111111111001110100",  "111111111001110011",  "111111111001110011",  "111111111001110010",  "111111111001110010",  "111111111001110010",  "111111111001110001",  "111111111001110001",  "111111111001110000",  "111111111001110000",  "111111111001101111",  "111111111001101111",  "111111111001101110",  "111111111001101110",  "111111111001101110",  "111111111001101101",  "111111111001101101",  "111111111001101100",  "111111111001101100",  "111111111001101011",  "111111111001101011",  "111111111001101011",  "111111111001101010",  "111111111001101010",  "111111111001101010",  "111111111001101001",  "111111111001101001",  "111111111001101000",  "111111111001101000",  "111111111001101000",  "111111111001100111",  "111111111001100111",  "111111111001100111",  "111111111001100110",  "111111111001100110",  "111111111001100110",  "111111111001100101",  "111111111001100101",  "111111111001100100",  "111111111001100100",  "111111111001100100",  "111111111001100100",  "111111111001100011",  "111111111001100011",  "111111111001100011",  "111111111001100010",  "111111111001100010",  "111111111001100010",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100000",  "111111111001100000",  "111111111001100000",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001010111",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011000",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011001",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011010",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011011",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011100",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011101",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011110",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001011111",  "111111111001100000",  "111111111001100000",  "111111111001100000",  "111111111001100000",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100001",  "111111111001100010",  "111111111001100010",  "111111111001100010",  "111111111001100011",  "111111111001100011",  "111111111001100011",  "111111111001100100",  "111111111001100100",  "111111111001100100",  "111111111001100101",  "111111111001100101",  "111111111001100101",  "111111111001100101",  "111111111001100110",  "111111111001100110",  "111111111001100110",  "111111111001100111",  "111111111001100111",  "111111111001101000",  "111111111001101000",  "111111111001101000",  "111111111001101001",  "111111111001101001",  "111111111001101001",  "111111111001101010",  "111111111001101010",  "111111111001101010",  "111111111001101011",  "111111111001101011",  "111111111001101100",  "111111111001101100",  "111111111001101100",  "111111111001101101",  "111111111001101101",  "111111111001101110",  "111111111001101110",  "111111111001101111",  "111111111001101111",  "111111111001101111",  "111111111001110000",  "111111111001110000",  "111111111001110001",  "111111111001110001",  "111111111001110010",  "111111111001110010",  "111111111001110010",  "111111111001110011",  "111111111001110011",  "111111111001110100",  "111111111001110100",  "111111111001110101",  "111111111001110101",  "111111111001110110",  "111111111001110110",  "111111111001110111",  "111111111001110111",  "111111111001111000",  "111111111001111000",  "111111111001111001",  "111111111001111001",  "111111111001111010",  "111111111001111010",  "111111111001111011",  "111111111001111011",  "111111111001111100",  "111111111001111100",  "111111111001111101",  "111111111001111101",  "111111111001111110",  "111111111001111110",  "111111111001111111",  "111111111001111111",  "111111111010000000",  "111111111010000000",  "111111111010000001",  "111111111010000010",  "111111111010000010",  "111111111010000011",  "111111111010000011",  "111111111010000100",  "111111111010000100",  "111111111010000101",  "111111111010000110",  "111111111010000110",  "111111111010000111",  "111111111010000111",  "111111111010001000",  "111111111010001000",  "111111111010001001",  "111111111010001010",  "111111111010001010",  "111111111010001011",  "111111111010001100",  "111111111010001100",  "111111111010001101",  "111111111010001101",  "111111111010001110",  "111111111010001111",  "111111111010001111",  "111111111010010000",  "111111111010010001",  "111111111010010001",  "111111111010010010",  "111111111010010010",  "111111111010010011",  "111111111010010100",  "111111111010010100",  "111111111010010101",  "111111111010010110",  "111111111010010110",  "111111111010010111",  "111111111010011000",  "111111111010011000",  "111111111010011001",  "111111111010011010",  "111111111010011010",  "111111111010011011",  "111111111010011100",  "111111111010011101",  "111111111010011101",  "111111111010011110",  "111111111010011111",  "111111111010011111",  "111111111010100000",  "111111111010100001",  "111111111010100001",  "111111111010100010",  "111111111010100011",  "111111111010100100",  "111111111010100100",  "111111111010100101",  "111111111010100110",  "111111111010100111",  "111111111010100111",  "111111111010101000",  "111111111010101001",  "111111111010101001",  "111111111010101010",  "111111111010101011",  "111111111010101100",  "111111111010101100",  "111111111010101101",  "111111111010101110",  "111111111010101111",  "111111111010110000",  "111111111010110000",  "111111111010110001",  "111111111010110010",  "111111111010110011",  "111111111010110011",  "111111111010110100",  "111111111010110101",  "111111111010110110",  "111111111010110111",  "111111111010110111",  "111111111010111000",  "111111111010111001",  "111111111010111010",  "111111111010111011",  "111111111010111011",  "111111111010111100",  "111111111010111101",  "111111111010111110",  "111111111010111111",  "111111111011000000",  "111111111011000000",  "111111111011000001",  "111111111011000010",  "111111111011000011",  "111111111011000100",  "111111111011000101",  "111111111011000101",  "111111111011000110",  "111111111011000111",  "111111111011001000",  "111111111011001001",  "111111111011001010",  "111111111011001010",  "111111111011001011",  "111111111011001100",  "111111111011001101",  "111111111011001110",  "111111111011001111",  "111111111011010000",  "111111111011010001",  "111111111011010001",  "111111111011010010",  "111111111011010011",  "111111111011010100",  "111111111011010101",  "111111111011010110",  "111111111011010111",  "111111111011011000",  "111111111011011001",  "111111111011011001",  "111111111011011010",  "111111111011011011",  "111111111011011100",  "111111111011011101",  "111111111011011110",  "111111111011011111",  "111111111011100000",  "111111111011100001",  "111111111011100010",  "111111111011100011",  "111111111011100011",  "111111111011100100",  "111111111011100101",  "111111111011100110",  "111111111011100111",  "111111111011101000",  "111111111011101001",  "111111111011101010",  "111111111011101011",  "111111111011101100",  "111111111011101101",  "111111111011101110",  "111111111011101111",  "111111111011110000",  "111111111011110001",  "111111111011110010",  "111111111011110011",  "111111111011110011",  "111111111011110100",  "111111111011110101",  "111111111011110110",  "111111111011110111",  "111111111011111000",  "111111111011111001",  "111111111011111010",  "111111111011111011",  "111111111011111100",  "111111111011111101",  "111111111011111110",  "111111111011111111",  "111111111100000000",  "111111111100000001",  "111111111100000010",  "111111111100000011",  "111111111100000100",  "111111111100000101",  "111111111100000110",  "111111111100000111",  "111111111100001000",  "111111111100001001",  "111111111100001010",  "111111111100001011",  "111111111100001100",  "111111111100001101",  "111111111100001110",  "111111111100001111",  "111111111100010000",  "111111111100010001",  "111111111100010010",  "111111111100010011",  "111111111100010100",  "111111111100010101",  "111111111100010110",  "111111111100010111",  "111111111100011000",  "111111111100011001",  "111111111100011011",  "111111111100011100",  "111111111100011101",  "111111111100011110",  "111111111100011111",  "111111111100100000",  "111111111100100001",  "111111111100100010",  "111111111100100011",  "111111111100100100",  "111111111100100101",  "111111111100100110",  "111111111100100111",  "111111111100101000",  "111111111100101001",  "111111111100101010",  "111111111100101011",  "111111111100101100",  "111111111100101101",  "111111111100101110",  "111111111100110000",  "111111111100110001",  "111111111100110010",  "111111111100110011",  "111111111100110100",  "111111111100110101",  "111111111100110110",  "111111111100110111",  "111111111100111000",  "111111111100111001",  "111111111100111010",  "111111111100111011",  "111111111100111100",  "111111111100111110",  "111111111100111111",  "111111111101000000",  "111111111101000001",  "111111111101000010",  "111111111101000011",  "111111111101000100",  "111111111101000101",  "111111111101000110",  "111111111101000111",  "111111111101001000",  "111111111101001010",  "111111111101001011",  "111111111101001100",  "111111111101001101",  "111111111101001110",  "111111111101001111",  "111111111101010000",  "111111111101010001",  "111111111101010010",  "111111111101010011",  "111111111101010101",  "111111111101010110",  "111111111101010111",  "111111111101011000",  "111111111101011001",  "111111111101011010",  "111111111101011011",  "111111111101011100",  "111111111101011110",  "111111111101011111",  "111111111101100000",  "111111111101100001",  "111111111101100010",  "111111111101100011",  "111111111101100100",  "111111111101100101",  "111111111101100110",  "111111111101101000",  "111111111101101001",  "111111111101101010",  "111111111101101011",  "111111111101101100",  "111111111101101101",  "111111111101101110",  "111111111101110000",  "111111111101110001",  "111111111101110010",  "111111111101110011",  "111111111101110100",  "111111111101110101",  "111111111101110110",  "111111111101110111",  "111111111101111001",  "111111111101111010",  "111111111101111011",  "111111111101111100",  "111111111101111101",  "111111111101111110",  "111111111101111111",  "111111111110000001",  "111111111110000010",  "111111111110000011",  "111111111110000100",  "111111111110000101",  "111111111110000110",  "111111111110001000",  "111111111110001001",  "111111111110001010",  "111111111110001011",  "111111111110001100",  "111111111110001101",  "111111111110001110",  "111111111110010000",  "111111111110010001",  "111111111110010010",  "111111111110010011",  "111111111110010100",  "111111111110010101",  "111111111110010110",  "111111111110011000",  "111111111110011001",  "111111111110011010",  "111111111110011011",  "111111111110011100",  "111111111110011101",  "111111111110011111",  "111111111110100000",  "111111111110100001",  "111111111110100010",  "111111111110100011",  "111111111110100100",  "111111111110100110",  "111111111110100111",  "111111111110101000",  "111111111110101001",  "111111111110101010",  "111111111110101011",  "111111111110101100",  "111111111110101110",  "111111111110101111",  "111111111110110000",  "111111111110110001",  "111111111110110010",  "111111111110110011",  "111111111110110101",  "111111111110110110",  "111111111110110111",  "111111111110111000",  "111111111110111001",  "111111111110111010",  "111111111110111100",  "111111111110111101",  "111111111110111110",  "111111111110111111",  "111111111111000000",  "111111111111000001",  "111111111111000011",  "111111111111000100",  "111111111111000101",  "111111111111000110",  "111111111111000111",  "111111111111001000",  "111111111111001010",  "111111111111001011",  "111111111111001100",  "111111111111001101",  "111111111111001110",  "111111111111001111",  "111111111111010001",  "111111111111010010",  "111111111111010011",  "111111111111010100",  "111111111111010101",  "111111111111010110",  "111111111111011000",  "111111111111011001",  "111111111111011010",  "111111111111011011",  "111111111111011100",  "111111111111011101",  "111111111111011110",  "111111111111100000",  "111111111111100001",  "111111111111100010",  "111111111111100011",  "111111111111100100",  "111111111111100101",  "111111111111100111",  "111111111111101000",  "111111111111101001",  "111111111111101010",  "111111111111101011",  "111111111111101100",  "111111111111101110",  "111111111111101111",  "111111111111110000",  "111111111111110001",  "111111111111110010",  "111111111111110011",  "111111111111110100",  "111111111111110110",  "111111111111110111",  "111111111111111000",  "111111111111111001",  "111111111111111010",  "111111111111111011",  "111111111111111101",  "111111111111111110",  "111111111111111111"),("000000000000000000",  "000000000000000001",  "000000000000000010",  "000000000000000011",  "000000000000000101",  "000000000000000110",  "000000000000000111",  "000000000000001000",  "000000000000001001",  "000000000000001010",  "000000000000001011",  "000000000000001101",  "000000000000001110",  "000000000000001111",  "000000000000010000",  "000000000000010001",  "000000000000010010",  "000000000000010011",  "000000000000010101",  "000000000000010110",  "000000000000010111",  "000000000000011000",  "000000000000011001",  "000000000000011010",  "000000000000011011",  "000000000000011101",  "000000000000011110",  "000000000000011111",  "000000000000100000",  "000000000000100001",  "000000000000100010",  "000000000000100011",  "000000000000100100",  "000000000000100110",  "000000000000100111",  "000000000000101000",  "000000000000101001",  "000000000000101010",  "000000000000101011",  "000000000000101100",  "000000000000101101",  "000000000000101111",  "000000000000110000",  "000000000000110001",  "000000000000110010",  "000000000000110011",  "000000000000110100",  "000000000000110101",  "000000000000110110",  "000000000000110111",  "000000000000111001",  "000000000000111010",  "000000000000111011",  "000000000000111100",  "000000000000111101",  "000000000000111110",  "000000000000111111",  "000000000001000000",  "000000000001000001",  "000000000001000010",  "000000000001000100",  "000000000001000101",  "000000000001000110",  "000000000001000111",  "000000000001001000",  "000000000001001001",  "000000000001001010",  "000000000001001011",  "000000000001001100",  "000000000001001101",  "000000000001001110",  "000000000001010000",  "000000000001010001",  "000000000001010010",  "000000000001010011",  "000000000001010100",  "000000000001010101",  "000000000001010110",  "000000000001010111",  "000000000001011000",  "000000000001011001",  "000000000001011010",  "000000000001011011",  "000000000001011100",  "000000000001011110",  "000000000001011111",  "000000000001100000",  "000000000001100001",  "000000000001100010",  "000000000001100011",  "000000000001100100",  "000000000001100101",  "000000000001100110",  "000000000001100111",  "000000000001101000",  "000000000001101001",  "000000000001101010",  "000000000001101011",  "000000000001101100",  "000000000001101101",  "000000000001101110",  "000000000001101111",  "000000000001110000",  "000000000001110001",  "000000000001110011",  "000000000001110100",  "000000000001110101",  "000000000001110110",  "000000000001110111",  "000000000001111000",  "000000000001111001",  "000000000001111010",  "000000000001111011",  "000000000001111100",  "000000000001111101",  "000000000001111110",  "000000000001111111",  "000000000010000000",  "000000000010000001",  "000000000010000010",  "000000000010000011",  "000000000010000100",  "000000000010000101",  "000000000010000110",  "000000000010000111",  "000000000010001000",  "000000000010001001",  "000000000010001010",  "000000000010001011",  "000000000010001100",  "000000000010001101",  "000000000010001110",  "000000000010001111",  "000000000010010000",  "000000000010010001",  "000000000010010010",  "000000000010010011",  "000000000010010100",  "000000000010010101",  "000000000010010110",  "000000000010010111",  "000000000010011000",  "000000000010011001",  "000000000010011010",  "000000000010011011",  "000000000010011100",  "000000000010011101",  "000000000010011101",  "000000000010011110",  "000000000010011111",  "000000000010100000",  "000000000010100001",  "000000000010100010",  "000000000010100011",  "000000000010100100",  "000000000010100101",  "000000000010100110",  "000000000010100111",  "000000000010101000",  "000000000010101001",  "000000000010101010",  "000000000010101011",  "000000000010101100",  "000000000010101101",  "000000000010101101",  "000000000010101110",  "000000000010101111",  "000000000010110000",  "000000000010110001",  "000000000010110010",  "000000000010110011",  "000000000010110100",  "000000000010110101",  "000000000010110110",  "000000000010110111",  "000000000010111000",  "000000000010111000",  "000000000010111001",  "000000000010111010",  "000000000010111011",  "000000000010111100",  "000000000010111101",  "000000000010111110",  "000000000010111111",  "000000000011000000",  "000000000011000000",  "000000000011000001",  "000000000011000010",  "000000000011000011",  "000000000011000100",  "000000000011000101",  "000000000011000110",  "000000000011000111",  "000000000011000111",  "000000000011001000",  "000000000011001001",  "000000000011001010",  "000000000011001011",  "000000000011001100",  "000000000011001100",  "000000000011001101",  "000000000011001110",  "000000000011001111",  "000000000011010000",  "000000000011010001",  "000000000011010010",  "000000000011010010",  "000000000011010011",  "000000000011010100",  "000000000011010101",  "000000000011010110",  "000000000011010110",  "000000000011010111",  "000000000011011000",  "000000000011011001",  "000000000011011010",  "000000000011011011",  "000000000011011011",  "000000000011011100",  "000000000011011101",  "000000000011011110",  "000000000011011111",  "000000000011011111",  "000000000011100000",  "000000000011100001",  "000000000011100010",  "000000000011100010",  "000000000011100011",  "000000000011100100",  "000000000011100101",  "000000000011100110",  "000000000011100110",  "000000000011100111",  "000000000011101000",  "000000000011101001",  "000000000011101001",  "000000000011101010",  "000000000011101011",  "000000000011101100",  "000000000011101100",  "000000000011101101",  "000000000011101110",  "000000000011101111",  "000000000011101111",  "000000000011110000",  "000000000011110001",  "000000000011110010",  "000000000011110010",  "000000000011110011",  "000000000011110100",  "000000000011110100",  "000000000011110101",  "000000000011110110",  "000000000011110111",  "000000000011110111",  "000000000011111000",  "000000000011111001",  "000000000011111001",  "000000000011111010",  "000000000011111011",  "000000000011111011",  "000000000011111100",  "000000000011111101",  "000000000011111110",  "000000000011111110",  "000000000011111111",  "000000000100000000",  "000000000100000000",  "000000000100000001",  "000000000100000010",  "000000000100000010",  "000000000100000011",  "000000000100000100",  "000000000100000100",  "000000000100000101",  "000000000100000110",  "000000000100000110",  "000000000100000111",  "000000000100000111",  "000000000100001000",  "000000000100001001",  "000000000100001001",  "000000000100001010",  "000000000100001011",  "000000000100001011",  "000000000100001100",  "000000000100001100",  "000000000100001101",  "000000000100001110",  "000000000100001110",  "000000000100001111",  "000000000100010000",  "000000000100010000",  "000000000100010001",  "000000000100010001",  "000000000100010010",  "000000000100010011",  "000000000100010011",  "000000000100010100",  "000000000100010100",  "000000000100010101",  "000000000100010101",  "000000000100010110",  "000000000100010111",  "000000000100010111",  "000000000100011000",  "000000000100011000",  "000000000100011001",  "000000000100011001",  "000000000100011010",  "000000000100011010",  "000000000100011011",  "000000000100011100",  "000000000100011100",  "000000000100011101",  "000000000100011101",  "000000000100011110",  "000000000100011110",  "000000000100011111",  "000000000100011111",  "000000000100100000",  "000000000100100000",  "000000000100100001",  "000000000100100001",  "000000000100100010",  "000000000100100010",  "000000000100100011",  "000000000100100011",  "000000000100100100",  "000000000100100100",  "000000000100100101",  "000000000100100101",  "000000000100100110",  "000000000100100110",  "000000000100100111",  "000000000100100111",  "000000000100101000",  "000000000100101000",  "000000000100101001",  "000000000100101001",  "000000000100101010",  "000000000100101010",  "000000000100101010",  "000000000100101011",  "000000000100101011",  "000000000100101100",  "000000000100101100",  "000000000100101101",  "000000000100101101",  "000000000100101110",  "000000000100101110",  "000000000100101110",  "000000000100101111",  "000000000100101111",  "000000000100110000",  "000000000100110000",  "000000000100110001",  "000000000100110001",  "000000000100110001",  "000000000100110010",  "000000000100110010",  "000000000100110011",  "000000000100110011",  "000000000100110011",  "000000000100110100",  "000000000100110100",  "000000000100110100",  "000000000100110101",  "000000000100110101",  "000000000100110110",  "000000000100110110",  "000000000100110110",  "000000000100110111",  "000000000100110111",  "000000000100110111",  "000000000100111000",  "000000000100111000",  "000000000100111000",  "000000000100111001",  "000000000100111001",  "000000000100111001",  "000000000100111010",  "000000000100111010",  "000000000100111010",  "000000000100111011",  "000000000100111011",  "000000000100111011",  "000000000100111100",  "000000000100111100",  "000000000100111100",  "000000000100111101",  "000000000100111101",  "000000000100111101",  "000000000100111101",  "000000000100111110",  "000000000100111110",  "000000000100111110",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000101000000",  "000000000101000000",  "000000000101000000",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001011",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001010",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001001",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101001000",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000111",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000110",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000101",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000100",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000011",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000010",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000001",  "000000000101000000",  "000000000101000000",  "000000000101000000",  "000000000101000000",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000100111111",  "000000000100111110",  "000000000100111110",  "000000000100111110",  "000000000100111110",  "000000000100111101",  "000000000100111101",  "000000000100111101",  "000000000100111100",  "000000000100111100",  "000000000100111100",  "000000000100111011",  "000000000100111011",  "000000000100111011",  "000000000100111011",  "000000000100111010",  "000000000100111010",  "000000000100111010",  "000000000100111001",  "000000000100111001",  "000000000100111001",  "000000000100111000",  "000000000100111000",  "000000000100111000",  "000000000100110111",  "000000000100110111",  "000000000100110111",  "000000000100110110",  "000000000100110110",  "000000000100110110",  "000000000100110101",  "000000000100110101",  "000000000100110100",  "000000000100110100",  "000000000100110100",  "000000000100110011",  "000000000100110011",  "000000000100110011",  "000000000100110010",  "000000000100110010",  "000000000100110010",  "000000000100110001",  "000000000100110001",  "000000000100110000",  "000000000100110000",  "000000000100110000",  "000000000100101111",  "000000000100101111",  "000000000100101110",  "000000000100101110",  "000000000100101110",  "000000000100101101",  "000000000100101101",  "000000000100101100",  "000000000100101100",  "000000000100101011",  "000000000100101011",  "000000000100101011",  "000000000100101010",  "000000000100101010",  "000000000100101001",  "000000000100101001",  "000000000100101000",  "000000000100101000",  "000000000100101000",  "000000000100100111",  "000000000100100111",  "000000000100100110",  "000000000100100110",  "000000000100100101",  "000000000100100101",  "000000000100100100",  "000000000100100100",  "000000000100100011",  "000000000100100011",  "000000000100100010",  "000000000100100010",  "000000000100100001",  "000000000100100001",  "000000000100100001",  "000000000100100000",  "000000000100100000",  "000000000100011111",  "000000000100011111",  "000000000100011110",  "000000000100011110",  "000000000100011101",  "000000000100011101",  "000000000100011100",  "000000000100011100",  "000000000100011011",  "000000000100011011",  "000000000100011010",  "000000000100011001",  "000000000100011001",  "000000000100011000",  "000000000100011000",  "000000000100010111",  "000000000100010111",  "000000000100010110",  "000000000100010110",  "000000000100010101",  "000000000100010101",  "000000000100010100",  "000000000100010100",  "000000000100010011",  "000000000100010011",  "000000000100010010",  "000000000100010001",  "000000000100010001",  "000000000100010000",  "000000000100010000",  "000000000100001111",  "000000000100001111",  "000000000100001110",  "000000000100001101",  "000000000100001101",  "000000000100001100",  "000000000100001100",  "000000000100001011",  "000000000100001011",  "000000000100001010",  "000000000100001001",  "000000000100001001",  "000000000100001000",  "000000000100001000",  "000000000100000111",  "000000000100000110",  "000000000100000110",  "000000000100000101",  "000000000100000101",  "000000000100000100",  "000000000100000011",  "000000000100000011",  "000000000100000010",  "000000000100000010",  "000000000100000001",  "000000000100000000",  "000000000100000000",  "000000000011111111",  "000000000011111111",  "000000000011111110",  "000000000011111101",  "000000000011111101",  "000000000011111100",  "000000000011111011",  "000000000011111011",  "000000000011111010",  "000000000011111001",  "000000000011111001",  "000000000011111000",  "000000000011111000",  "000000000011110111",  "000000000011110110",  "000000000011110110",  "000000000011110101",  "000000000011110100",  "000000000011110100",  "000000000011110011",  "000000000011110010",  "000000000011110010",  "000000000011110001",  "000000000011110000",  "000000000011110000",  "000000000011101111",  "000000000011101110",  "000000000011101110",  "000000000011101101",  "000000000011101100",  "000000000011101100",  "000000000011101011",  "000000000011101010",  "000000000011101001",  "000000000011101001",  "000000000011101000",  "000000000011100111",  "000000000011100111",  "000000000011100110",  "000000000011100101",  "000000000011100101",  "000000000011100100",  "000000000011100011",  "000000000011100010",  "000000000011100010",  "000000000011100001",  "000000000011100000",  "000000000011100000",  "000000000011011111",  "000000000011011110",  "000000000011011101",  "000000000011011101",  "000000000011011100",  "000000000011011011",  "000000000011011011",  "000000000011011010",  "000000000011011001",  "000000000011011000",  "000000000011011000",  "000000000011010111",  "000000000011010110",  "000000000011010101",  "000000000011010101",  "000000000011010100",  "000000000011010011",  "000000000011010010",  "000000000011010010",  "000000000011010001",  "000000000011010000",  "000000000011010000",  "000000000011001111",  "000000000011001110",  "000000000011001101",  "000000000011001100",  "000000000011001100",  "000000000011001011",  "000000000011001010",  "000000000011001001",  "000000000011001001",  "000000000011001000",  "000000000011000111",  "000000000011000110",  "000000000011000110",  "000000000011000101",  "000000000011000100",  "000000000011000011",  "000000000011000011",  "000000000011000010",  "000000000011000001",  "000000000011000000",  "000000000010111111",  "000000000010111111",  "000000000010111110",  "000000000010111101",  "000000000010111100",  "000000000010111011",  "000000000010111011",  "000000000010111010",  "000000000010111001",  "000000000010111000",  "000000000010110111",  "000000000010110111",  "000000000010110110",  "000000000010110101",  "000000000010110100",  "000000000010110011",  "000000000010110011",  "000000000010110010",  "000000000010110001",  "000000000010110000",  "000000000010101111",  "000000000010101111",  "000000000010101110",  "000000000010101101",  "000000000010101100",  "000000000010101011",  "000000000010101011",  "000000000010101010",  "000000000010101001",  "000000000010101000",  "000000000010100111",  "000000000010100110",  "000000000010100110",  "000000000010100101",  "000000000010100100",  "000000000010100011",  "000000000010100010",  "000000000010100010",  "000000000010100001",  "000000000010100000",  "000000000010011111",  "000000000010011110",  "000000000010011101",  "000000000010011101",  "000000000010011100",  "000000000010011011",  "000000000010011010",  "000000000010011001",  "000000000010011000",  "000000000010010111",  "000000000010010111",  "000000000010010110",  "000000000010010101",  "000000000010010100",  "000000000010010011",  "000000000010010010",  "000000000010010010",  "000000000010010001",  "000000000010010000",  "000000000010001111",  "000000000010001110",  "000000000010001101",  "000000000010001100",  "000000000010001100",  "000000000010001011",  "000000000010001010",  "000000000010001001",  "000000000010001000",  "000000000010000111",  "000000000010000110",  "000000000010000110",  "000000000010000101",  "000000000010000100",  "000000000010000011",  "000000000010000010",  "000000000010000001",  "000000000010000000",  "000000000010000000",  "000000000001111111",  "000000000001111110",  "000000000001111101",  "000000000001111100",  "000000000001111011",  "000000000001111010",  "000000000001111001",  "000000000001111001",  "000000000001111000",  "000000000001110111",  "000000000001110110",  "000000000001110101",  "000000000001110100",  "000000000001110011",  "000000000001110010",  "000000000001110010",  "000000000001110001",  "000000000001110000",  "000000000001101111",  "000000000001101110",  "000000000001101101",  "000000000001101100",  "000000000001101011",  "000000000001101011",  "000000000001101010",  "000000000001101001",  "000000000001101000",  "000000000001100111",  "000000000001100110",  "000000000001100101",  "000000000001100100",  "000000000001100011",  "000000000001100011",  "000000000001100010",  "000000000001100001",  "000000000001100000",  "000000000001011111",  "000000000001011110",  "000000000001011101",  "000000000001011100",  "000000000001011011",  "000000000001011011",  "000000000001011010",  "000000000001011001",  "000000000001011000",  "000000000001010111",  "000000000001010110",  "000000000001010101",  "000000000001010100",  "000000000001010011",  "000000000001010011",  "000000000001010010",  "000000000001010001",  "000000000001010000",  "000000000001001111",  "000000000001001110",  "000000000001001101",  "000000000001001100",  "000000000001001011",  "000000000001001010",  "000000000001001010",  "000000000001001001",  "000000000001001000",  "000000000001000111",  "000000000001000110",  "000000000001000101",  "000000000001000100",  "000000000001000011",  "000000000001000010",  "000000000001000001",  "000000000001000001",  "000000000001000000",  "000000000000111111",  "000000000000111110",  "000000000000111101",  "000000000000111100",  "000000000000111011",  "000000000000111010",  "000000000000111001",  "000000000000111000",  "000000000000111000",  "000000000000110111",  "000000000000110110",  "000000000000110101",  "000000000000110100",  "000000000000110011",  "000000000000110010",  "000000000000110001",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101101",  "000000000000101100",  "000000000000101011",  "000000000000101010",  "000000000000101001",  "000000000000101000",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100100",  "000000000000100011",  "000000000000100010",  "000000000000100001",  "000000000000100000",  "000000000000011111",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011011",  "000000000000011010",  "000000000000011001",  "000000000000011000",  "000000000000010111",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010011",  "000000000000010010",  "000000000000010001",  "000000000000010000",  "000000000000001111",  "000000000000001110",  "000000000000001101",  "000000000000001100",  "000000000000001100",  "000000000000001011",  "000000000000001010",  "000000000000001001",  "000000000000001000",  "000000000000000111",  "000000000000000110",  "000000000000000101",  "000000000000000100",  "000000000000000100",  "000000000000000011",  "000000000000000010",  "000000000000000001"),("000000000000000000",  "111111111111111111",  "111111111111111110",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111010",  "111111111111111001",  "111111111111111000",  "111111111111110111",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110011",  "111111111111110010",  "111111111111110001",  "111111111111110000",  "111111111111101111",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101011",  "111111111111101010",  "111111111111101001",  "111111111111101000",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100100",  "111111111111100011",  "111111111111100010",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011110",  "111111111111011101",  "111111111111011100",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011000",  "111111111111010111",  "111111111111010110",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010010",  "111111111111010001",  "111111111111010000",  "111111111111001111",  "111111111111001110",  "111111111111001110",  "111111111111001101",  "111111111111001100",  "111111111111001011",  "111111111111001010",  "111111111111001001",  "111111111111001000",  "111111111111001000",  "111111111111000111",  "111111111111000110",  "111111111111000101",  "111111111111000100",  "111111111111000011",  "111111111111000011",  "111111111111000010",  "111111111111000001",  "111111111111000000",  "111111111110111111",  "111111111110111110",  "111111111110111110",  "111111111110111101",  "111111111110111100",  "111111111110111011",  "111111111110111010",  "111111111110111001",  "111111111110111001",  "111111111110111000",  "111111111110110111",  "111111111110110110",  "111111111110110101",  "111111111110110101",  "111111111110110100",  "111111111110110011",  "111111111110110010",  "111111111110110001",  "111111111110110001",  "111111111110110000",  "111111111110101111",  "111111111110101110",  "111111111110101101",  "111111111110101100",  "111111111110101100",  "111111111110101011",  "111111111110101010",  "111111111110101001",  "111111111110101000",  "111111111110101000",  "111111111110100111",  "111111111110100110",  "111111111110100101",  "111111111110100100",  "111111111110100100",  "111111111110100011",  "111111111110100010",  "111111111110100001",  "111111111110100001",  "111111111110100000",  "111111111110011111",  "111111111110011110",  "111111111110011101",  "111111111110011101",  "111111111110011100",  "111111111110011011",  "111111111110011010",  "111111111110011010",  "111111111110011001",  "111111111110011000",  "111111111110010111",  "111111111110010110",  "111111111110010110",  "111111111110010101",  "111111111110010100",  "111111111110010011",  "111111111110010011",  "111111111110010010",  "111111111110010001",  "111111111110010000",  "111111111110010000",  "111111111110001111",  "111111111110001110",  "111111111110001101",  "111111111110001101",  "111111111110001100",  "111111111110001011",  "111111111110001010",  "111111111110001010",  "111111111110001001",  "111111111110001000",  "111111111110000111",  "111111111110000111",  "111111111110000110",  "111111111110000101",  "111111111110000100",  "111111111110000100",  "111111111110000011",  "111111111110000010",  "111111111110000010",  "111111111110000001",  "111111111110000000",  "111111111101111111",  "111111111101111111",  "111111111101111110",  "111111111101111101",  "111111111101111100",  "111111111101111100",  "111111111101111011",  "111111111101111010",  "111111111101111010",  "111111111101111001",  "111111111101111000",  "111111111101111000",  "111111111101110111",  "111111111101110110",  "111111111101110101",  "111111111101110101",  "111111111101110100",  "111111111101110011",  "111111111101110011",  "111111111101110010",  "111111111101110001",  "111111111101110001",  "111111111101110000",  "111111111101101111",  "111111111101101111",  "111111111101101110",  "111111111101101101",  "111111111101101100",  "111111111101101100",  "111111111101101011",  "111111111101101010",  "111111111101101010",  "111111111101101001",  "111111111101101000",  "111111111101101000",  "111111111101100111",  "111111111101100110",  "111111111101100110",  "111111111101100101",  "111111111101100100",  "111111111101100100",  "111111111101100011",  "111111111101100011",  "111111111101100010",  "111111111101100001",  "111111111101100001",  "111111111101100000",  "111111111101011111",  "111111111101011111",  "111111111101011110",  "111111111101011101",  "111111111101011101",  "111111111101011100",  "111111111101011100",  "111111111101011011",  "111111111101011010",  "111111111101011010",  "111111111101011001",  "111111111101011000",  "111111111101011000",  "111111111101010111",  "111111111101010111",  "111111111101010110",  "111111111101010101",  "111111111101010101",  "111111111101010100",  "111111111101010100",  "111111111101010011",  "111111111101010010",  "111111111101010010",  "111111111101010001",  "111111111101010001",  "111111111101010000",  "111111111101001111",  "111111111101001111",  "111111111101001110",  "111111111101001110",  "111111111101001101",  "111111111101001100",  "111111111101001100",  "111111111101001011",  "111111111101001011",  "111111111101001010",  "111111111101001010",  "111111111101001001",  "111111111101001000",  "111111111101001000",  "111111111101000111",  "111111111101000111",  "111111111101000110",  "111111111101000110",  "111111111101000101",  "111111111101000100",  "111111111101000100",  "111111111101000011",  "111111111101000011",  "111111111101000010",  "111111111101000010",  "111111111101000001",  "111111111101000001",  "111111111101000000",  "111111111101000000",  "111111111100111111",  "111111111100111111",  "111111111100111110",  "111111111100111110",  "111111111100111101",  "111111111100111100",  "111111111100111100",  "111111111100111011",  "111111111100111011",  "111111111100111010",  "111111111100111010",  "111111111100111001",  "111111111100111001",  "111111111100111000",  "111111111100111000",  "111111111100110111",  "111111111100110111",  "111111111100110110",  "111111111100110110",  "111111111100110101",  "111111111100110101",  "111111111100110100",  "111111111100110100",  "111111111100110011",  "111111111100110011",  "111111111100110011",  "111111111100110010",  "111111111100110010",  "111111111100110001",  "111111111100110001",  "111111111100110000",  "111111111100110000",  "111111111100101111",  "111111111100101111",  "111111111100101110",  "111111111100101110",  "111111111100101101",  "111111111100101101",  "111111111100101101",  "111111111100101100",  "111111111100101100",  "111111111100101011",  "111111111100101011",  "111111111100101010",  "111111111100101010",  "111111111100101001",  "111111111100101001",  "111111111100101001",  "111111111100101000",  "111111111100101000",  "111111111100100111",  "111111111100100111",  "111111111100100110",  "111111111100100110",  "111111111100100110",  "111111111100100101",  "111111111100100101",  "111111111100100100",  "111111111100100100",  "111111111100100100",  "111111111100100011",  "111111111100100011",  "111111111100100010",  "111111111100100010",  "111111111100100010",  "111111111100100001",  "111111111100100001",  "111111111100100000",  "111111111100100000",  "111111111100100000",  "111111111100011111",  "111111111100011111",  "111111111100011111",  "111111111100011110",  "111111111100011110",  "111111111100011110",  "111111111100011101",  "111111111100011101",  "111111111100011100",  "111111111100011100",  "111111111100011100",  "111111111100011011",  "111111111100011011",  "111111111100011011",  "111111111100011010",  "111111111100011010",  "111111111100011010",  "111111111100011001",  "111111111100011001",  "111111111100011001",  "111111111100011000",  "111111111100011000",  "111111111100011000",  "111111111100010111",  "111111111100010111",  "111111111100010111",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010101",  "111111111100010101",  "111111111100010101",  "111111111100010100",  "111111111100010100",  "111111111100010100",  "111111111100010011",  "111111111100010011",  "111111111100010011",  "111111111100010011",  "111111111100010010",  "111111111100010010",  "111111111100010010",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000010",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000011",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000100",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000101",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000110",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100000111",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001000",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001001",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001010",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001011",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001100",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001101",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001110",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100001111",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100010000",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010001",  "111111111100010010",  "111111111100010010",  "111111111100010010",  "111111111100010010",  "111111111100010011",  "111111111100010011",  "111111111100010011",  "111111111100010100",  "111111111100010100",  "111111111100010100",  "111111111100010100",  "111111111100010101",  "111111111100010101",  "111111111100010101",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010110",  "111111111100010111",  "111111111100010111",  "111111111100010111",  "111111111100011000",  "111111111100011000",  "111111111100011000",  "111111111100011001",  "111111111100011001",  "111111111100011001",  "111111111100011001",  "111111111100011010",  "111111111100011010",  "111111111100011010",  "111111111100011011",  "111111111100011011",  "111111111100011011",  "111111111100011100",  "111111111100011100",  "111111111100011100",  "111111111100011101",  "111111111100011101",  "111111111100011101",  "111111111100011110",  "111111111100011110",  "111111111100011110",  "111111111100011111",  "111111111100011111",  "111111111100100000",  "111111111100100000",  "111111111100100000",  "111111111100100001",  "111111111100100001",  "111111111100100001",  "111111111100100010",  "111111111100100010",  "111111111100100010",  "111111111100100011",  "111111111100100011",  "111111111100100100",  "111111111100100100",  "111111111100100100",  "111111111100100101",  "111111111100100101",  "111111111100100101",  "111111111100100110",  "111111111100100110",  "111111111100100111",  "111111111100100111",  "111111111100100111",  "111111111100101000",  "111111111100101000",  "111111111100101001",  "111111111100101001",  "111111111100101001",  "111111111100101010",  "111111111100101010",  "111111111100101011",  "111111111100101011",  "111111111100101011",  "111111111100101100",  "111111111100101100",  "111111111100101101",  "111111111100101101",  "111111111100101101",  "111111111100101110",  "111111111100101110",  "111111111100101111",  "111111111100101111",  "111111111100110000",  "111111111100110000",  "111111111100110000",  "111111111100110001",  "111111111100110001",  "111111111100110010",  "111111111100110010",  "111111111100110011",  "111111111100110011",  "111111111100110100",  "111111111100110100",  "111111111100110100",  "111111111100110101",  "111111111100110101",  "111111111100110110",  "111111111100110110",  "111111111100110111",  "111111111100110111",  "111111111100111000",  "111111111100111000",  "111111111100111001",  "111111111100111001",  "111111111100111001",  "111111111100111010",  "111111111100111010",  "111111111100111011",  "111111111100111011",  "111111111100111100",  "111111111100111100",  "111111111100111101",  "111111111100111101",  "111111111100111110",  "111111111100111110",  "111111111100111111",  "111111111100111111",  "111111111101000000",  "111111111101000000",  "111111111101000001",  "111111111101000001",  "111111111101000010",  "111111111101000010",  "111111111101000011",  "111111111101000011",  "111111111101000100",  "111111111101000100",  "111111111101000101",  "111111111101000101",  "111111111101000110",  "111111111101000110",  "111111111101000111",  "111111111101000111",  "111111111101001000",  "111111111101001000",  "111111111101001001",  "111111111101001001",  "111111111101001010",  "111111111101001010",  "111111111101001011",  "111111111101001011",  "111111111101001100",  "111111111101001100",  "111111111101001101",  "111111111101001101",  "111111111101001110",  "111111111101001110",  "111111111101001111",  "111111111101001111",  "111111111101010000",  "111111111101010001",  "111111111101010001",  "111111111101010010",  "111111111101010010",  "111111111101010011",  "111111111101010011",  "111111111101010100",  "111111111101010100",  "111111111101010101",  "111111111101010101",  "111111111101010110",  "111111111101010111",  "111111111101010111",  "111111111101011000",  "111111111101011000",  "111111111101011001",  "111111111101011001",  "111111111101011010",  "111111111101011010",  "111111111101011011",  "111111111101011100",  "111111111101011100",  "111111111101011101",  "111111111101011101",  "111111111101011110",  "111111111101011110",  "111111111101011111",  "111111111101100000",  "111111111101100000",  "111111111101100001",  "111111111101100001",  "111111111101100010",  "111111111101100010",  "111111111101100011",  "111111111101100100",  "111111111101100100",  "111111111101100101",  "111111111101100101",  "111111111101100110",  "111111111101100110",  "111111111101100111",  "111111111101101000",  "111111111101101000",  "111111111101101001",  "111111111101101001",  "111111111101101010",  "111111111101101011",  "111111111101101011",  "111111111101101100",  "111111111101101100",  "111111111101101101",  "111111111101101110",  "111111111101101110",  "111111111101101111",  "111111111101101111",  "111111111101110000",  "111111111101110001",  "111111111101110001",  "111111111101110010",  "111111111101110010",  "111111111101110011",  "111111111101110100",  "111111111101110100",  "111111111101110101",  "111111111101110101",  "111111111101110110",  "111111111101110111",  "111111111101110111",  "111111111101111000",  "111111111101111000",  "111111111101111001",  "111111111101111010",  "111111111101111010",  "111111111101111011",  "111111111101111100",  "111111111101111100",  "111111111101111101",  "111111111101111101",  "111111111101111110",  "111111111101111111",  "111111111101111111",  "111111111110000000",  "111111111110000001",  "111111111110000001",  "111111111110000010",  "111111111110000010",  "111111111110000011",  "111111111110000100",  "111111111110000100",  "111111111110000101",  "111111111110000110",  "111111111110000110",  "111111111110000111",  "111111111110001000",  "111111111110001000",  "111111111110001001",  "111111111110001001",  "111111111110001010",  "111111111110001011",  "111111111110001011",  "111111111110001100",  "111111111110001101",  "111111111110001101",  "111111111110001110",  "111111111110001111",  "111111111110001111",  "111111111110010000",  "111111111110010001",  "111111111110010001",  "111111111110010010",  "111111111110010010",  "111111111110010011",  "111111111110010100",  "111111111110010100",  "111111111110010101",  "111111111110010110",  "111111111110010110",  "111111111110010111",  "111111111110011000",  "111111111110011000",  "111111111110011001",  "111111111110011010",  "111111111110011010",  "111111111110011011",  "111111111110011100",  "111111111110011100",  "111111111110011101",  "111111111110011110",  "111111111110011110",  "111111111110011111",  "111111111110100000",  "111111111110100000",  "111111111110100001",  "111111111110100010",  "111111111110100010",  "111111111110100011",  "111111111110100100",  "111111111110100100",  "111111111110100101",  "111111111110100110",  "111111111110100110",  "111111111110100111",  "111111111110101000",  "111111111110101000",  "111111111110101001",  "111111111110101010",  "111111111110101010",  "111111111110101011",  "111111111110101100",  "111111111110101100",  "111111111110101101",  "111111111110101110",  "111111111110101110",  "111111111110101111",  "111111111110110000",  "111111111110110000",  "111111111110110001",  "111111111110110010",  "111111111110110010",  "111111111110110011",  "111111111110110100",  "111111111110110100",  "111111111110110101",  "111111111110110110",  "111111111110110110",  "111111111110110111",  "111111111110111000",  "111111111110111000",  "111111111110111001",  "111111111110111010",  "111111111110111010",  "111111111110111011",  "111111111110111100",  "111111111110111100",  "111111111110111101",  "111111111110111110",  "111111111110111111",  "111111111110111111",  "111111111111000000",  "111111111111000001",  "111111111111000001",  "111111111111000010",  "111111111111000011",  "111111111111000011",  "111111111111000100",  "111111111111000101",  "111111111111000101",  "111111111111000110",  "111111111111000111",  "111111111111000111",  "111111111111001000",  "111111111111001001",  "111111111111001001",  "111111111111001010",  "111111111111001011",  "111111111111001011",  "111111111111001100",  "111111111111001101",  "111111111111001110",  "111111111111001110",  "111111111111001111",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111111",  "111111111111111111"),("000000000000000000",  "000000000000000001",  "000000000000000001",  "000000000000000010",  "000000000000000011",  "000000000000000011",  "000000000000000100",  "000000000000000101",  "000000000000000101",  "000000000000000110",  "000000000000000111",  "000000000000000111",  "000000000000001000",  "000000000000001001",  "000000000000001001",  "000000000000001010",  "000000000000001011",  "000000000000001011",  "000000000000001100",  "000000000000001101",  "000000000000001101",  "000000000000001110",  "000000000000001111",  "000000000000001111",  "000000000000010000",  "000000000000010001",  "000000000000010001",  "000000000000010010",  "000000000000010011",  "000000000000010011",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010111",  "000000000000010111",  "000000000000011000",  "000000000000011001",  "000000000000011001",  "000000000000011010",  "000000000000011011",  "000000000000011011",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011111",  "000000000000011111",  "000000000000100000",  "000000000000100000",  "000000000000100001",  "000000000000100010",  "000000000000100010",  "000000000000100011",  "000000000000100100",  "000000000000100100",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000101000",  "000000000000101000",  "000000000000101001",  "000000000000101001",  "000000000000101010",  "000000000000101011",  "000000000000101011",  "000000000000101100",  "000000000000101101",  "000000000000101101",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110000",  "000000000000110001",  "000000000000110010",  "000000000000110010",  "000000000000110011",  "000000000000110100",  "000000000000110100",  "000000000000110101",  "000000000000110101",  "000000000000110110",  "000000000000110111",  "000000000000110111",  "000000000000111000",  "000000000000111001",  "000000000000111001",  "000000000000111010",  "000000000000111010",  "000000000000111011",  "000000000000111100",  "000000000000111100",  "000000000000111101",  "000000000000111101",  "000000000000111110",  "000000000000111111",  "000000000000111111",  "000000000001000000",  "000000000001000001",  "000000000001000001",  "000000000001000010",  "000000000001000010",  "000000000001000011",  "000000000001000100",  "000000000001000100",  "000000000001000101",  "000000000001000101",  "000000000001000110",  "000000000001000111",  "000000000001000111",  "000000000001001000",  "000000000001001000",  "000000000001001001",  "000000000001001010",  "000000000001001010",  "000000000001001011",  "000000000001001011",  "000000000001001100",  "000000000001001100",  "000000000001001101",  "000000000001001110",  "000000000001001110",  "000000000001001111",  "000000000001001111",  "000000000001010000",  "000000000001010001",  "000000000001010001",  "000000000001010010",  "000000000001010010",  "000000000001010011",  "000000000001010011",  "000000000001010100",  "000000000001010101",  "000000000001010101",  "000000000001010110",  "000000000001010110",  "000000000001010111",  "000000000001010111",  "000000000001011000",  "000000000001011001",  "000000000001011001",  "000000000001011010",  "000000000001011010",  "000000000001011011",  "000000000001011011",  "000000000001011100",  "000000000001011100",  "000000000001011101",  "000000000001011110",  "000000000001011110",  "000000000001011111",  "000000000001011111",  "000000000001100000",  "000000000001100000",  "000000000001100001",  "000000000001100001",  "000000000001100010",  "000000000001100010",  "000000000001100011",  "000000000001100100",  "000000000001100100",  "000000000001100101",  "000000000001100101",  "000000000001100110",  "000000000001100110",  "000000000001100111",  "000000000001100111",  "000000000001101000",  "000000000001101000",  "000000000001101001",  "000000000001101001",  "000000000001101010",  "000000000001101010",  "000000000001101011",  "000000000001101011",  "000000000001101100",  "000000000001101101",  "000000000001101101",  "000000000001101110",  "000000000001101110",  "000000000001101111",  "000000000001101111",  "000000000001110000",  "000000000001110000",  "000000000001110001",  "000000000001110001",  "000000000001110010",  "000000000001110010",  "000000000001110011",  "000000000001110011",  "000000000001110100",  "000000000001110100",  "000000000001110101",  "000000000001110101",  "000000000001110110",  "000000000001110110",  "000000000001110111",  "000000000001110111",  "000000000001111000",  "000000000001111000",  "000000000001111001",  "000000000001111001",  "000000000001111010",  "000000000001111010",  "000000000001111010",  "000000000001111011",  "000000000001111011",  "000000000001111100",  "000000000001111100",  "000000000001111101",  "000000000001111101",  "000000000001111110",  "000000000001111110",  "000000000001111111",  "000000000001111111",  "000000000010000000",  "000000000010000000",  "000000000010000001",  "000000000010000001",  "000000000010000010",  "000000000010000010",  "000000000010000010",  "000000000010000011",  "000000000010000011",  "000000000010000100",  "000000000010000100",  "000000000010000101",  "000000000010000101",  "000000000010000110",  "000000000010000110",  "000000000010000110",  "000000000010000111",  "000000000010000111",  "000000000010001000",  "000000000010001000",  "000000000010001001",  "000000000010001001",  "000000000010001001",  "000000000010001010",  "000000000010001010",  "000000000010001011",  "000000000010001011",  "000000000010001100",  "000000000010001100",  "000000000010001100",  "000000000010001101",  "000000000010001101",  "000000000010001110",  "000000000010001110",  "000000000010001111",  "000000000010001111",  "000000000010001111",  "000000000010010000",  "000000000010010000",  "000000000010010001",  "000000000010010001",  "000000000010010001",  "000000000010010010",  "000000000010010010",  "000000000010010011",  "000000000010010011",  "000000000010010011",  "000000000010010100",  "000000000010010100",  "000000000010010101",  "000000000010010101",  "000000000010010101",  "000000000010010110",  "000000000010010110",  "000000000010010110",  "000000000010010111",  "000000000010010111",  "000000000010011000",  "000000000010011000",  "000000000010011000",  "000000000010011001",  "000000000010011001",  "000000000010011001",  "000000000010011010",  "000000000010011010",  "000000000010011010",  "000000000010011011",  "000000000010011011",  "000000000010011100",  "000000000010011100",  "000000000010011100",  "000000000010011101",  "000000000010011101",  "000000000010011101",  "000000000010011110",  "000000000010011110",  "000000000010011110",  "000000000010011111",  "000000000010011111",  "000000000010011111",  "000000000010100000",  "000000000010100000",  "000000000010100000",  "000000000010100001",  "000000000010100001",  "000000000010100001",  "000000000010100010",  "000000000010100010",  "000000000010100010",  "000000000010100011",  "000000000010100011",  "000000000010100011",  "000000000010100100",  "000000000010100100",  "000000000010100100",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100110",  "000000000010100110",  "000000000010100110",  "000000000010100111",  "000000000010100111",  "000000000010100111",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010101001",  "000000000010101001",  "000000000010101001",  "000000000010101010",  "000000000010101010",  "000000000010101010",  "000000000010101010",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111111",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111110",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111101",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111100",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111011",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111010",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111001",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010111000",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110111",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110110",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110101",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110100",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110011",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110010",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110001",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010110000",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010101111",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101110",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101101",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101100",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101011",  "000000000010101010",  "000000000010101010",  "000000000010101010",  "000000000010101001",  "000000000010101001",  "000000000010101001",  "000000000010101001",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010101000",  "000000000010100111",  "000000000010100111",  "000000000010100111",  "000000000010100111",  "000000000010100110",  "000000000010100110",  "000000000010100110",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100101",  "000000000010100100",  "000000000010100100",  "000000000010100100",  "000000000010100011",  "000000000010100011",  "000000000010100011",  "000000000010100010",  "000000000010100010",  "000000000010100010",  "000000000010100010",  "000000000010100001",  "000000000010100001",  "000000000010100001",  "000000000010100000",  "000000000010100000",  "000000000010100000",  "000000000010011111",  "000000000010011111",  "000000000010011111",  "000000000010011110",  "000000000010011110",  "000000000010011110",  "000000000010011110",  "000000000010011101",  "000000000010011101",  "000000000010011101",  "000000000010011100",  "000000000010011100",  "000000000010011100",  "000000000010011011",  "000000000010011011",  "000000000010011011",  "000000000010011010",  "000000000010011010",  "000000000010011010",  "000000000010011001",  "000000000010011001",  "000000000010011001",  "000000000010011000",  "000000000010011000",  "000000000010011000",  "000000000010010111",  "000000000010010111",  "000000000010010111",  "000000000010010110",  "000000000010010110",  "000000000010010101",  "000000000010010101",  "000000000010010101",  "000000000010010100",  "000000000010010100",  "000000000010010100",  "000000000010010011",  "000000000010010011",  "000000000010010011",  "000000000010010010",  "000000000010010010",  "000000000010010010",  "000000000010010001",  "000000000010010001",  "000000000010010000",  "000000000010010000",  "000000000010010000",  "000000000010001111",  "000000000010001111",  "000000000010001111",  "000000000010001110",  "000000000010001110",  "000000000010001110",  "000000000010001101",  "000000000010001101",  "000000000010001100",  "000000000010001100",  "000000000010001100",  "000000000010001011",  "000000000010001011",  "000000000010001010",  "000000000010001010",  "000000000010001010",  "000000000010001001",  "000000000010001001",  "000000000010001001",  "000000000010001000",  "000000000010001000",  "000000000010000111",  "000000000010000111",  "000000000010000111",  "000000000010000110",  "000000000010000110",  "000000000010000101",  "000000000010000101",  "000000000010000101",  "000000000010000100",  "000000000010000100",  "000000000010000011",  "000000000010000011",  "000000000010000011",  "000000000010000010",  "000000000010000010",  "000000000010000001",  "000000000010000001",  "000000000010000001",  "000000000010000000",  "000000000010000000",  "000000000001111111",  "000000000001111111",  "000000000001111110",  "000000000001111110",  "000000000001111110",  "000000000001111101",  "000000000001111101",  "000000000001111100",  "000000000001111100",  "000000000001111100",  "000000000001111011",  "000000000001111011",  "000000000001111010",  "000000000001111010",  "000000000001111001",  "000000000001111001",  "000000000001111001",  "000000000001111000",  "000000000001111000",  "000000000001110111",  "000000000001110111",  "000000000001110110",  "000000000001110110",  "000000000001110110",  "000000000001110101",  "000000000001110101",  "000000000001110100",  "000000000001110100",  "000000000001110011",  "000000000001110011",  "000000000001110010",  "000000000001110010",  "000000000001110010",  "000000000001110001",  "000000000001110001",  "000000000001110000",  "000000000001110000",  "000000000001101111",  "000000000001101111",  "000000000001101110",  "000000000001101110",  "000000000001101110",  "000000000001101101",  "000000000001101101",  "000000000001101100",  "000000000001101100",  "000000000001101011",  "000000000001101011",  "000000000001101010",  "000000000001101010",  "000000000001101001",  "000000000001101001",  "000000000001101001",  "000000000001101000",  "000000000001101000",  "000000000001100111",  "000000000001100111",  "000000000001100110",  "000000000001100110",  "000000000001100101",  "000000000001100101",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100011",  "000000000001100011",  "000000000001100010",  "000000000001100010",  "000000000001100001",  "000000000001100001",  "000000000001100000",  "000000000001100000",  "000000000001011111",  "000000000001011111",  "000000000001011110",  "000000000001011110",  "000000000001011101",  "000000000001011101",  "000000000001011100",  "000000000001011100",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011010",  "000000000001011010",  "000000000001011001",  "000000000001011001",  "000000000001011000",  "000000000001011000",  "000000000001010111",  "000000000001010111",  "000000000001010110",  "000000000001010110",  "000000000001010101",  "000000000001010101",  "000000000001010100",  "000000000001010100",  "000000000001010011",  "000000000001010011",  "000000000001010010",  "000000000001010010",  "000000000001010001",  "000000000001010001",  "000000000001010000",  "000000000001010000",  "000000000001001111",  "000000000001001111",  "000000000001001110",  "000000000001001110",  "000000000001001101",  "000000000001001101",  "000000000001001100",  "000000000001001100",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001010",  "000000000001001010",  "000000000001001001",  "000000000001001001",  "000000000001001000",  "000000000001001000",  "000000000001000111",  "000000000001000111",  "000000000001000110",  "000000000001000110",  "000000000001000101",  "000000000001000101",  "000000000001000100",  "000000000001000100",  "000000000001000011",  "000000000001000011",  "000000000001000010",  "000000000001000010",  "000000000001000001",  "000000000001000001",  "000000000001000000",  "000000000001000000",  "000000000000111111",  "000000000000111111",  "000000000000111110",  "000000000000111110",  "000000000000111101",  "000000000000111101",  "000000000000111100",  "000000000000111100",  "000000000000111011",  "000000000000111011",  "000000000000111010",  "000000000000111010",  "000000000000111001",  "000000000000111000",  "000000000000111000",  "000000000000110111",  "000000000000110111",  "000000000000110110",  "000000000000110110",  "000000000000110101",  "000000000000110101",  "000000000000110100",  "000000000000110100",  "000000000000110011",  "000000000000110011",  "000000000000110010",  "000000000000110010",  "000000000000110001",  "000000000000110001",  "000000000000110000",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101110",  "000000000000101101",  "000000000000101101",  "000000000000101100",  "000000000000101100",  "000000000000101011",  "000000000000101011",  "000000000000101010",  "000000000000101010",  "000000000000101001",  "000000000000101001",  "000000000000101000",  "000000000000101000",  "000000000000100111",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100101",  "000000000000100100",  "000000000000100100",  "000000000000100011",  "000000000000100011",  "000000000000100010",  "000000000000100010",  "000000000000100001",  "000000000000100001",  "000000000000100000",  "000000000000100000",  "000000000000011111",  "000000000000011110",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011100",  "000000000000011011",  "000000000000011011",  "000000000000011010",  "000000000000011010",  "000000000000011001",  "000000000000011001",  "000000000000011000",  "000000000000011000",  "000000000000010111",  "000000000000010111",  "000000000000010110",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010100",  "000000000000010011",  "000000000000010011",  "000000000000010010",  "000000000000010010",  "000000000000010001",  "000000000000010001",  "000000000000010000",  "000000000000010000",  "000000000000001111",  "000000000000001111",  "000000000000001110",  "000000000000001110",  "000000000000001101",  "000000000000001101",  "000000000000001100",  "000000000000001100",  "000000000000001011",  "000000000000001011",  "000000000000001010",  "000000000000001010",  "000000000000001001",  "000000000000001001",  "000000000000001000",  "000000000000001000",  "000000000000000111",  "000000000000000111",  "000000000000000110",  "000000000000000110",  "000000000000000101",  "000000000000000101",  "000000000000000100",  "000000000000000100",  "000000000000000011",  "000000000000000011",  "000000000000000010",  "000000000000000010",  "000000000000000001",  "000000000000000001"),("000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111001111",  "111111111111001111",  "111111111111001110",  "111111111111001110",  "111111111111001101",  "111111111111001101",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001011",  "111111111111001011",  "111111111111001010",  "111111111111001010",  "111111111111001001",  "111111111111001001",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111000111",  "111111111111000111",  "111111111111000110",  "111111111111000110",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000100",  "111111111111000100",  "111111111111000011",  "111111111111000011",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000001",  "111111111111000001",  "111111111111000000",  "111111111111000000",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111110",  "111111111110111110",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111100",  "111111111110111100",  "111111111110111011",  "111111111110111011",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111001",  "111111111110111001",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110110111",  "111111111110110111",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110101",  "111111111110110101",  "111111111110110100",  "111111111110110100",  "111111111110110100",  "111111111110110011",  "111111111110110011",  "111111111110110010",  "111111111110110010",  "111111111110110010",  "111111111110110001",  "111111111110110001",  "111111111110110001",  "111111111110110000",  "111111111110110000",  "111111111110101111",  "111111111110101111",  "111111111110101111",  "111111111110101110",  "111111111110101110",  "111111111110101101",  "111111111110101101",  "111111111110101101",  "111111111110101100",  "111111111110101100",  "111111111110101100",  "111111111110101011",  "111111111110101011",  "111111111110101010",  "111111111110101010",  "111111111110101010",  "111111111110101001",  "111111111110101001",  "111111111110101001",  "111111111110101000",  "111111111110101000",  "111111111110101000",  "111111111110100111",  "111111111110100111",  "111111111110100110",  "111111111110100110",  "111111111110100110",  "111111111110100101",  "111111111110100101",  "111111111110100101",  "111111111110100100",  "111111111110100100",  "111111111110100100",  "111111111110100011",  "111111111110100011",  "111111111110100011",  "111111111110100010",  "111111111110100010",  "111111111110100010",  "111111111110100001",  "111111111110100001",  "111111111110100001",  "111111111110100000",  "111111111110100000",  "111111111110100000",  "111111111110011111",  "111111111110011111",  "111111111110011111",  "111111111110011110",  "111111111110011110",  "111111111110011110",  "111111111110011101",  "111111111110011101",  "111111111110011101",  "111111111110011100",  "111111111110011100",  "111111111110011100",  "111111111110011011",  "111111111110011011",  "111111111110011011",  "111111111110011010",  "111111111110011010",  "111111111110011010",  "111111111110011001",  "111111111110011001",  "111111111110011001",  "111111111110011000",  "111111111110011000",  "111111111110011000",  "111111111110010111",  "111111111110010111",  "111111111110010111",  "111111111110010111",  "111111111110010110",  "111111111110010110",  "111111111110010110",  "111111111110010101",  "111111111110010101",  "111111111110010101",  "111111111110010100",  "111111111110010100",  "111111111110010100",  "111111111110010100",  "111111111110010011",  "111111111110010011",  "111111111110010011",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010001",  "111111111110010001",  "111111111110010001",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110001110",  "111111111110001110",  "111111111110001110",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110011",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110100",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110101",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110110",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101110111",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111000",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111001",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111010",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111011",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111100",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111101",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111110",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111101111111",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000000",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000001",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000010",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000011",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000100",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000101",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000110",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110000111",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001000",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001001",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001010",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001011",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001100",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001101",  "111111111110001110",  "111111111110001110",  "111111111110001110",  "111111111110001110",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110001111",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110010000",  "111111111110010001",  "111111111110010001",  "111111111110010001",  "111111111110010001",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010010",  "111111111110010011",  "111111111110010011",  "111111111110010011",  "111111111110010011",  "111111111110010100",  "111111111110010100",  "111111111110010100",  "111111111110010101",  "111111111110010101",  "111111111110010101",  "111111111110010101",  "111111111110010110",  "111111111110010110",  "111111111110010110",  "111111111110010110",  "111111111110010111",  "111111111110010111",  "111111111110010111",  "111111111110011000",  "111111111110011000",  "111111111110011000",  "111111111110011000",  "111111111110011001",  "111111111110011001",  "111111111110011001",  "111111111110011001",  "111111111110011010",  "111111111110011010",  "111111111110011010",  "111111111110011011",  "111111111110011011",  "111111111110011011",  "111111111110011011",  "111111111110011100",  "111111111110011100",  "111111111110011100",  "111111111110011101",  "111111111110011101",  "111111111110011101",  "111111111110011110",  "111111111110011110",  "111111111110011110",  "111111111110011110",  "111111111110011111",  "111111111110011111",  "111111111110011111",  "111111111110100000",  "111111111110100000",  "111111111110100000",  "111111111110100001",  "111111111110100001",  "111111111110100001",  "111111111110100001",  "111111111110100010",  "111111111110100010",  "111111111110100010",  "111111111110100011",  "111111111110100011",  "111111111110100011",  "111111111110100100",  "111111111110100100",  "111111111110100100",  "111111111110100100",  "111111111110100101",  "111111111110100101",  "111111111110100101",  "111111111110100110",  "111111111110100110",  "111111111110100110",  "111111111110100111",  "111111111110100111",  "111111111110100111",  "111111111110101000",  "111111111110101000",  "111111111110101000",  "111111111110101001",  "111111111110101001",  "111111111110101001",  "111111111110101010",  "111111111110101010",  "111111111110101010",  "111111111110101011",  "111111111110101011",  "111111111110101011",  "111111111110101011",  "111111111110101100",  "111111111110101100",  "111111111110101100",  "111111111110101101",  "111111111110101101",  "111111111110101101",  "111111111110101110",  "111111111110101110",  "111111111110101110",  "111111111110101111",  "111111111110101111",  "111111111110101111",  "111111111110110000",  "111111111110110000",  "111111111110110000",  "111111111110110001",  "111111111110110001",  "111111111110110001",  "111111111110110010",  "111111111110110010",  "111111111110110010",  "111111111110110011",  "111111111110110011",  "111111111110110011",  "111111111110110100",  "111111111110110100",  "111111111110110100",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110110",  "111111111110110110",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111110",  "111111111110111110",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000100",  "111111111111000100",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111001000",  "111111111111001000",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001100",  "111111111111001100",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111110",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000010",  "000000000000000010",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000110",  "000000000000000110",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001010",  "000000000000001010",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001110",  "000000000000001110",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010100",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111011",  "000000000000111011",  "000000000000111011",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111110",  "000000000000111110",  "000000000000111110",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100111",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100110",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100101",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100100",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100011",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100010",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100001",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001100000",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011111",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011110",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011101",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011100",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011011",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011010",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011001",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001011000",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010111",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010110",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010101",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010100",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010011",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010010",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010001",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001010000",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001111",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001110",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001101",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001100",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001011",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001010",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001001",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001001000",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001000111",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000110",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000101",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000100",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000011",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000010",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000001",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000001000000",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111111",  "000000000000111110",  "000000000000111110",  "000000000000111110",  "000000000000111110",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111101",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111100",  "000000000000111011",  "000000000000111011",  "000000000000111011",  "000000000000111011",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111010",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110101",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110110",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110110111",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111000",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111001",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111010",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111011",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111100",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111101",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111110",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111110111111",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000000",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000001",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000010",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000011",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000100",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000101",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000110",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111000111",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001000",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001001",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001010",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001011",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001100",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001101",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001110",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111001111",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "000000000000000000",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "000000000000000000",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111001",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000111000",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110111",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110110",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110101",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110100",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110011",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110010",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110001",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000110000",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101111",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101110",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101101",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101100",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101011",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101010",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101001",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000101000",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100111",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100110",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100101",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100100",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100011",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100010",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100001",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000100000",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011111",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011110",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011101",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011100",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011011",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011010",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011001",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000011000",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010111",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010110",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010101",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010100",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010011",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010010",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010001",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000010000",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001111",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001110",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001101",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001100",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001011",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001010",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001001",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000001000",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000111",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000110",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000101",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000100",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000011",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000010",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000001",  "000000000000000000",  "000000000000000000",  "000000000000000000"),("000000000000000000",  "000000000000000000",  "000000000000000000",  "000000000000000000",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010000",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010001",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010010",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010011",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010100",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010101",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010110",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111010111",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011000",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011001",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011010",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011011",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011100",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011101",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011110",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111011111",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100000",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100001",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100010",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100011",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100100",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100101",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100110",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111100111",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101000",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101001",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101010",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101011",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101100",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101101",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101110",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111101111",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110000",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110001",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110010",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110011",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110100",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110101",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110110",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111110111",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111000",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111001",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111010",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111011",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111100",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111101",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111110",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "111111111111111111",  "000000000000000000",  "000000000000000000",  "000000000000000000") );

end CoeffConstants;

package body CoeffConstants is
end CoeffConstants;
